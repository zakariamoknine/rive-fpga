// Generator : SpinalHDL dev    git head : 84ef7b5b6278854e0e80738536f72c64fa14b730
// Component : VexiiRiscv
// Git hash  : fc927f9311a0f0710a1a90b88b62d9d5a020e9c6

`timescale 1ns/1ps

module VexiiRiscv (
  output wire          LsuL1Axi4Plugin_logic_axi_aw_valid,
  input  wire          LsuL1Axi4Plugin_logic_axi_aw_ready,
  output wire [31:0]   LsuL1Axi4Plugin_logic_axi_aw_payload_addr,
  output wire [7:0]    LsuL1Axi4Plugin_logic_axi_aw_payload_len,
  output wire [2:0]    LsuL1Axi4Plugin_logic_axi_aw_payload_size,
  output wire [1:0]    LsuL1Axi4Plugin_logic_axi_aw_payload_burst,
  output wire [3:0]    LsuL1Axi4Plugin_logic_axi_aw_payload_cache,
  output wire [2:0]    LsuL1Axi4Plugin_logic_axi_aw_payload_prot,
  output wire          LsuL1Axi4Plugin_logic_axi_w_valid,
  input  wire          LsuL1Axi4Plugin_logic_axi_w_ready,
  output wire [63:0]   LsuL1Axi4Plugin_logic_axi_w_payload_data,
  output wire [7:0]    LsuL1Axi4Plugin_logic_axi_w_payload_strb,
  output wire          LsuL1Axi4Plugin_logic_axi_w_payload_last,
  input  wire          LsuL1Axi4Plugin_logic_axi_b_valid,
  output wire          LsuL1Axi4Plugin_logic_axi_b_ready,
  input  wire [1:0]    LsuL1Axi4Plugin_logic_axi_b_payload_resp,
  output wire          LsuL1Axi4Plugin_logic_axi_ar_valid,
  input  wire          LsuL1Axi4Plugin_logic_axi_ar_ready,
  output wire [31:0]   LsuL1Axi4Plugin_logic_axi_ar_payload_addr,
  output wire [7:0]    LsuL1Axi4Plugin_logic_axi_ar_payload_len,
  output wire [2:0]    LsuL1Axi4Plugin_logic_axi_ar_payload_size,
  output wire [1:0]    LsuL1Axi4Plugin_logic_axi_ar_payload_burst,
  output wire [3:0]    LsuL1Axi4Plugin_logic_axi_ar_payload_cache,
  output wire [2:0]    LsuL1Axi4Plugin_logic_axi_ar_payload_prot,
  input  wire          LsuL1Axi4Plugin_logic_axi_r_valid,
  output wire          LsuL1Axi4Plugin_logic_axi_r_ready,
  input  wire [63:0]   LsuL1Axi4Plugin_logic_axi_r_payload_data,
  input  wire [1:0]    LsuL1Axi4Plugin_logic_axi_r_payload_resp,
  input  wire          LsuL1Axi4Plugin_logic_axi_r_payload_last,
  input  wire [63:0]   PrivilegedPlugin_logic_rdtime,
  input  wire          PrivilegedPlugin_logic_harts_0_int_m_timer /* verilator public */ ,
  input  wire          PrivilegedPlugin_logic_harts_0_int_m_software /* verilator public */ ,
  input  wire          PrivilegedPlugin_logic_harts_0_int_m_external /* verilator public */ ,
  input  wire          PrivilegedPlugin_logic_harts_0_int_s_external /* verilator public */ ,
  output wire          FetchL1Axi4Plugin_logic_axi_ar_valid,
  input  wire          FetchL1Axi4Plugin_logic_axi_ar_ready,
  output wire [31:0]   FetchL1Axi4Plugin_logic_axi_ar_payload_addr,
  output wire [7:0]    FetchL1Axi4Plugin_logic_axi_ar_payload_len,
  output wire [2:0]    FetchL1Axi4Plugin_logic_axi_ar_payload_size,
  output wire [1:0]    FetchL1Axi4Plugin_logic_axi_ar_payload_burst,
  output wire [3:0]    FetchL1Axi4Plugin_logic_axi_ar_payload_cache,
  output wire [2:0]    FetchL1Axi4Plugin_logic_axi_ar_payload_prot,
  input  wire          FetchL1Axi4Plugin_logic_axi_r_valid,
  output wire          FetchL1Axi4Plugin_logic_axi_r_ready,
  input  wire [63:0]   FetchL1Axi4Plugin_logic_axi_r_payload_data,
  input  wire [1:0]    FetchL1Axi4Plugin_logic_axi_r_payload_resp,
  input  wire          FetchL1Axi4Plugin_logic_axi_r_payload_last,
  output wire          LsuCachelessAxi4Plugin_logic_axi_aw_valid,
  input  wire          LsuCachelessAxi4Plugin_logic_axi_aw_ready,
  output wire [31:0]   LsuCachelessAxi4Plugin_logic_axi_aw_payload_addr,
  output wire [2:0]    LsuCachelessAxi4Plugin_logic_axi_aw_payload_size,
  output wire [3:0]    LsuCachelessAxi4Plugin_logic_axi_aw_payload_cache,
  output wire [2:0]    LsuCachelessAxi4Plugin_logic_axi_aw_payload_prot,
  output wire          LsuCachelessAxi4Plugin_logic_axi_w_valid,
  input  wire          LsuCachelessAxi4Plugin_logic_axi_w_ready,
  output wire [63:0]   LsuCachelessAxi4Plugin_logic_axi_w_payload_data,
  output wire [7:0]    LsuCachelessAxi4Plugin_logic_axi_w_payload_strb,
  output wire          LsuCachelessAxi4Plugin_logic_axi_w_payload_last,
  input  wire          LsuCachelessAxi4Plugin_logic_axi_b_valid,
  output wire          LsuCachelessAxi4Plugin_logic_axi_b_ready,
  input  wire [1:0]    LsuCachelessAxi4Plugin_logic_axi_b_payload_resp,
  output wire          LsuCachelessAxi4Plugin_logic_axi_ar_valid,
  input  wire          LsuCachelessAxi4Plugin_logic_axi_ar_ready,
  output wire [31:0]   LsuCachelessAxi4Plugin_logic_axi_ar_payload_addr,
  output wire [2:0]    LsuCachelessAxi4Plugin_logic_axi_ar_payload_size,
  output wire [3:0]    LsuCachelessAxi4Plugin_logic_axi_ar_payload_cache,
  output wire [2:0]    LsuCachelessAxi4Plugin_logic_axi_ar_payload_prot,
  input  wire          LsuCachelessAxi4Plugin_logic_axi_r_valid,
  output wire          LsuCachelessAxi4Plugin_logic_axi_r_ready,
  input  wire [63:0]   LsuCachelessAxi4Plugin_logic_axi_r_payload_data,
  input  wire [1:0]    LsuCachelessAxi4Plugin_logic_axi_r_payload_resp,
  input  wire          LsuCachelessAxi4Plugin_logic_axi_r_payload_last,
  input  wire          clk,
  input  wire          reset
);
  localparam EnvPluginOp_ECALL = 3'd0;
  localparam EnvPluginOp_EBREAK = 3'd1;
  localparam EnvPluginOp_PRIV_RET = 3'd2;
  localparam EnvPluginOp_FENCE_I = 3'd3;
  localparam EnvPluginOp_SFENCE_VMA = 3'd4;
  localparam EnvPluginOp_WFI = 3'd5;
  localparam BranchPlugin_BranchCtrlEnum_B = 2'd0;
  localparam BranchPlugin_BranchCtrlEnum_JAL = 2'd1;
  localparam BranchPlugin_BranchCtrlEnum_JALR = 2'd2;
  localparam IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 = 2'd0;
  localparam IntAluPlugin_AluBitwiseCtrlEnum_OR_1 = 2'd1;
  localparam IntAluPlugin_AluBitwiseCtrlEnum_AND_1 = 2'd2;
  localparam IntAluPlugin_AluBitwiseCtrlEnum_ZERO = 2'd3;
  localparam LsuL1CmdOpcode_LSU = 3'd0;
  localparam LsuL1CmdOpcode_ACCESS_1 = 3'd1;
  localparam LsuL1CmdOpcode_STORE_BUFFER = 3'd2;
  localparam LsuL1CmdOpcode_FLUSH = 3'd3;
  localparam LsuL1CmdOpcode_PREFETCH = 3'd4;
  localparam LsuPlugin_logic_flusher_IDLE = 2'd0;
  localparam LsuPlugin_logic_flusher_CMD = 2'd1;
  localparam LsuPlugin_logic_flusher_COMPLETION = 2'd2;
  localparam TrapPlugin_logic_harts_0_trap_fsm_RESET = 4'd0;
  localparam TrapPlugin_logic_harts_0_trap_fsm_RUNNING = 4'd1;
  localparam TrapPlugin_logic_harts_0_trap_fsm_COMPUTE = 4'd2;
  localparam TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC = 4'd3;
  localparam TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL = 4'd4;
  localparam TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC = 4'd5;
  localparam TrapPlugin_logic_harts_0_trap_fsm_TRAP_WAIT = 4'd6;
  localparam TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY = 4'd7;
  localparam TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC = 4'd8;
  localparam TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY = 4'd9;
  localparam TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP = 4'd10;
  localparam TrapPlugin_logic_harts_0_trap_fsm_JUMP = 4'd11;
  localparam TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH = 4'd12;
  localparam TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH = 4'd13;
  localparam MmuPlugin_logic_refill_BOOT = 4'd0;
  localparam MmuPlugin_logic_refill_IDLE = 4'd1;
  localparam MmuPlugin_logic_refill_CMD_0 = 4'd2;
  localparam MmuPlugin_logic_refill_CMD_1 = 4'd3;
  localparam MmuPlugin_logic_refill_CMD_2 = 4'd4;
  localparam MmuPlugin_logic_refill_RSP_0 = 4'd5;
  localparam MmuPlugin_logic_refill_RSP_1 = 4'd6;
  localparam MmuPlugin_logic_refill_RSP_2 = 4'd7;
  localparam MmuPlugin_logic_refill_DONE_0 = 4'd8;
  localparam MmuPlugin_logic_refill_DONE_1 = 4'd9;
  localparam MmuPlugin_logic_refill_DONE_2 = 4'd10;
  localparam CsrAccessPlugin_logic_fsm_IDLE = 2'd0;
  localparam CsrAccessPlugin_logic_fsm_READ = 2'd1;
  localparam CsrAccessPlugin_logic_fsm_WRITE = 2'd2;
  localparam CsrAccessPlugin_logic_fsm_COMPLETION = 2'd3;
  localparam PerformanceCounterPlugin_logic_fsm_BOOT = 3'd0;
  localparam PerformanceCounterPlugin_logic_fsm_IDLE = 3'd1;
  localparam PerformanceCounterPlugin_logic_fsm_READ_LOW = 3'd2;
  localparam PerformanceCounterPlugin_logic_fsm_CALC_LOW = 3'd3;
  localparam PerformanceCounterPlugin_logic_fsm_CSR_WRITE = 3'd4;

  reg                 early0_DivPlugin_logic_processing_div_io_cmd_valid;
  reg                 LsuPlugin_logic_flusher_arbiter_io_output_ready;
  wire                LsuPlugin_logic_onAddress0_arbiter_io_output_ready;
  reg                 MmuPlugin_logic_refill_arbiter_io_output_ready;
  reg                 MmuPlugin_logic_invalidate_arbiter_io_output_ready;
  reg                 integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_valid;
  reg        [4:0]    integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_address;
  reg        [63:0]   integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_data;
  wire       [37:0]   BtbPlugin_logic_ras_mem_stack_spinal_port0;
  reg        [63:0]   LsuL1Plugin_logic_banks_0_mem_spinal_port1;
  reg        [63:0]   LsuL1Plugin_logic_banks_1_mem_spinal_port1;
  reg        [21:0]   LsuL1Plugin_logic_ways_0_mem_spinal_port1;
  reg        [21:0]   LsuL1Plugin_logic_ways_1_mem_spinal_port1;
  reg        [2:0]    LsuL1Plugin_logic_shared_mem_spinal_port1;
  reg        [63:0]   LsuL1Plugin_logic_writeback_victimBuffer_spinal_port1;
  reg        [63:0]   FetchL1Plugin_logic_banks_0_mem_spinal_port1;
  reg        [63:0]   FetchL1Plugin_logic_banks_1_mem_spinal_port1;
  reg        [21:0]   FetchL1Plugin_logic_ways_0_mem_spinal_port1;
  reg        [21:0]   FetchL1Plugin_logic_ways_1_mem_spinal_port1;
  reg        [0:0]    FetchL1Plugin_logic_plru_mem_spinal_port1;
  reg        [3:0]    GSharePlugin_logic_mem_banks_0_spinal_port1;
  reg        [57:0]   BtbPlugin_logic_mem_spinal_port1;
  wire       [46:0]   FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_0_spinal_port1;
  wire       [46:0]   FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_1_spinal_port1;
  wire       [28:0]   FetchL1Plugin_logic_translationStorage_logic_sl_1_ways_0_spinal_port1;
  wire       [46:0]   LsuPlugin_logic_translationStorage_logic_sl_0_ways_0_spinal_port1;
  wire       [46:0]   LsuPlugin_logic_translationStorage_logic_sl_0_ways_1_spinal_port1;
  wire       [46:0]   LsuPlugin_logic_translationStorage_logic_sl_0_ways_2_spinal_port1;
  wire       [28:0]   LsuPlugin_logic_translationStorage_logic_sl_1_ways_0_spinal_port1;
  reg        [63:0]   CsrRamPlugin_logic_mem_spinal_port1;
  wire                early0_DivPlugin_logic_processing_div_io_cmd_ready;
  wire                early0_DivPlugin_logic_processing_div_io_rsp_valid;
  wire       [63:0]   early0_DivPlugin_logic_processing_div_io_rsp_payload_result;
  wire       [63:0]   early0_DivPlugin_logic_processing_div_io_rsp_payload_remain;
  wire                LsuPlugin_logic_flusher_arbiter_io_inputs_0_ready;
  wire                LsuPlugin_logic_flusher_arbiter_io_output_valid;
  wire       [0:0]    LsuPlugin_logic_flusher_arbiter_io_chosenOH;
  wire                LsuPlugin_logic_onAddress0_arbiter_io_inputs_0_ready;
  wire                LsuPlugin_logic_onAddress0_arbiter_io_inputs_1_ready;
  wire                LsuPlugin_logic_onAddress0_arbiter_io_inputs_2_ready;
  wire                LsuPlugin_logic_onAddress0_arbiter_io_output_valid;
  wire       [2:0]    LsuPlugin_logic_onAddress0_arbiter_io_output_payload_op;
  wire       [38:0]   LsuPlugin_logic_onAddress0_arbiter_io_output_payload_address;
  wire       [1:0]    LsuPlugin_logic_onAddress0_arbiter_io_output_payload_size;
  wire                LsuPlugin_logic_onAddress0_arbiter_io_output_payload_load;
  wire                LsuPlugin_logic_onAddress0_arbiter_io_output_payload_store;
  wire                LsuPlugin_logic_onAddress0_arbiter_io_output_payload_atomic;
  wire                LsuPlugin_logic_onAddress0_arbiter_io_output_payload_clean;
  wire                LsuPlugin_logic_onAddress0_arbiter_io_output_payload_invalidate;
  wire       [11:0]   LsuPlugin_logic_onAddress0_arbiter_io_output_payload_storeId;
  wire       [1:0]    LsuPlugin_logic_onAddress0_arbiter_io_chosen;
  wire       [2:0]    LsuPlugin_logic_onAddress0_arbiter_io_chosenOH;
  wire                streamArbiter_5_io_inputs_0_ready;
  wire                streamArbiter_5_io_output_valid;
  wire       [38:0]   streamArbiter_5_io_output_payload_pcOnLastSlice;
  wire       [38:0]   streamArbiter_5_io_output_payload_pcTarget;
  wire                streamArbiter_5_io_output_payload_taken;
  wire                streamArbiter_5_io_output_payload_isBranch;
  wire                streamArbiter_5_io_output_payload_isPush;
  wire                streamArbiter_5_io_output_payload_isPop;
  wire                streamArbiter_5_io_output_payload_wasWrong;
  wire                streamArbiter_5_io_output_payload_badPredictedTarget;
  wire       [11:0]   streamArbiter_5_io_output_payload_history;
  wire       [15:0]   streamArbiter_5_io_output_payload_uopId;
  wire       [1:0]    streamArbiter_5_io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    streamArbiter_5_io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  wire       [0:0]    streamArbiter_5_io_chosenOH;
  wire                MmuPlugin_logic_refill_arbiter_io_inputs_0_ready;
  wire                MmuPlugin_logic_refill_arbiter_io_output_valid;
  wire       [38:0]   MmuPlugin_logic_refill_arbiter_io_output_payload_address;
  wire       [0:0]    MmuPlugin_logic_refill_arbiter_io_output_payload_storageId;
  wire                MmuPlugin_logic_refill_arbiter_io_output_payload_storageEnable;
  wire       [0:0]    MmuPlugin_logic_refill_arbiter_io_chosenOH;
  wire                MmuPlugin_logic_invalidate_arbiter_io_inputs_0_ready;
  wire                MmuPlugin_logic_invalidate_arbiter_io_output_valid;
  wire       [0:0]    MmuPlugin_logic_invalidate_arbiter_io_chosenOH;
  wire       [63:0]   integer_RegFilePlugin_logic_regfile_fpga_io_reads_0_data;
  wire       [63:0]   integer_RegFilePlugin_logic_regfile_fpga_io_reads_1_data;
  wire       [20:0]   _zz_PmpPlugin_logic_entries_0_napot_24;
  wire       [20:0]   _zz_PmpPlugin_logic_entries_1_napot_24;
  wire       [20:0]   _zz_PmpPlugin_logic_entries_2_napot_24;
  wire       [20:0]   _zz_PmpPlugin_logic_entries_3_napot_24;
  wire       [63:0]   _zz_early0_IntAluPlugin_logic_alu_result;
  wire       [63:0]   _zz_early0_IntAluPlugin_logic_alu_result_1;
  wire       [63:0]   _zz_early0_IntAluPlugin_logic_alu_result_2;
  wire       [63:0]   _zz_early0_IntAluPlugin_logic_alu_result_3;
  wire       [63:0]   _zz_early0_IntAluPlugin_logic_alu_result_4;
  wire       [0:0]    _zz_early0_IntAluPlugin_logic_alu_result_5;
  wire       [5:0]    _zz_early0_BarrelShifterPlugin_logic_shift_amplitude;
  wire       [63:0]   _zz_early0_BarrelShifterPlugin_logic_shift_reversed;
  wire                _zz_early0_BarrelShifterPlugin_logic_shift_reversed_1;
  wire       [0:0]    _zz_early0_BarrelShifterPlugin_logic_shift_reversed_2;
  wire       [52:0]   _zz_early0_BarrelShifterPlugin_logic_shift_reversed_3;
  wire                _zz_early0_BarrelShifterPlugin_logic_shift_reversed_4;
  wire       [0:0]    _zz_early0_BarrelShifterPlugin_logic_shift_reversed_5;
  wire       [41:0]   _zz_early0_BarrelShifterPlugin_logic_shift_reversed_6;
  wire                _zz_early0_BarrelShifterPlugin_logic_shift_reversed_7;
  wire       [0:0]    _zz_early0_BarrelShifterPlugin_logic_shift_reversed_8;
  wire       [30:0]   _zz_early0_BarrelShifterPlugin_logic_shift_reversed_9;
  wire                _zz_early0_BarrelShifterPlugin_logic_shift_reversed_10;
  wire       [0:0]    _zz_early0_BarrelShifterPlugin_logic_shift_reversed_11;
  wire       [19:0]   _zz_early0_BarrelShifterPlugin_logic_shift_reversed_12;
  wire                _zz_early0_BarrelShifterPlugin_logic_shift_reversed_13;
  wire       [0:0]    _zz_early0_BarrelShifterPlugin_logic_shift_reversed_14;
  wire       [8:0]    _zz_early0_BarrelShifterPlugin_logic_shift_reversed_15;
  wire       [64:0]   _zz_early0_BarrelShifterPlugin_logic_shift_shifted;
  wire       [64:0]   _zz_early0_BarrelShifterPlugin_logic_shift_shifted_1;
  wire       [63:0]   _zz_early0_BarrelShifterPlugin_logic_shift_patched;
  wire                _zz_early0_BarrelShifterPlugin_logic_shift_patched_1;
  wire       [0:0]    _zz_early0_BarrelShifterPlugin_logic_shift_patched_2;
  wire       [52:0]   _zz_early0_BarrelShifterPlugin_logic_shift_patched_3;
  wire                _zz_early0_BarrelShifterPlugin_logic_shift_patched_4;
  wire       [0:0]    _zz_early0_BarrelShifterPlugin_logic_shift_patched_5;
  wire       [41:0]   _zz_early0_BarrelShifterPlugin_logic_shift_patched_6;
  wire                _zz_early0_BarrelShifterPlugin_logic_shift_patched_7;
  wire       [0:0]    _zz_early0_BarrelShifterPlugin_logic_shift_patched_8;
  wire       [30:0]   _zz_early0_BarrelShifterPlugin_logic_shift_patched_9;
  wire                _zz_early0_BarrelShifterPlugin_logic_shift_patched_10;
  wire       [0:0]    _zz_early0_BarrelShifterPlugin_logic_shift_patched_11;
  wire       [19:0]   _zz_early0_BarrelShifterPlugin_logic_shift_patched_12;
  wire                _zz_early0_BarrelShifterPlugin_logic_shift_patched_13;
  wire       [0:0]    _zz_early0_BarrelShifterPlugin_logic_shift_patched_14;
  wire       [8:0]    _zz_early0_BarrelShifterPlugin_logic_shift_patched_15;
  wire       [21:0]   _zz_LsuL1Plugin_logic_ways_0_mem_port;
  wire                _zz_LsuL1Plugin_logic_ways_0_mem_port_1;
  wire       [21:0]   _zz_LsuL1Plugin_logic_ways_1_mem_port;
  wire                _zz_LsuL1Plugin_logic_ways_1_mem_port_1;
  wire       [2:0]    _zz_LsuL1Plugin_logic_shared_mem_port;
  wire       [0:0]    _zz_LsuL1Plugin_logic_shared_lsuRead_rsp_plru_0_1;
  wire       [2:0]    _zz_LsuL1Plugin_logic_writeback_read_wordIndex;
  wire       [0:0]    _zz_LsuL1Plugin_logic_writeback_read_wordIndex_1;
  reg        [63:0]   _zz_LsuL1Plugin_logic_writeback_read_readedData;
  wire       [2:0]    _zz_LsuL1Plugin_logic_writeback_victimBuffer_port;
  wire       [2:0]    _zz_LsuL1Plugin_logic_writeback_write_wordIndex;
  wire       [0:0]    _zz_LsuL1Plugin_logic_writeback_write_wordIndex_1;
  wire       [1:0]    _zz_LsuL1Plugin_logic_lsu_ctrl_refillWayNeedWriteback;
  wire       [0:0]    _zz_LsuL1Plugin_logic_lsu_ctrl_doWrite;
  reg        [1:0]    _zz_56;
  wire       [1:0]    _zz_57;
  reg        [1:0]    _zz_58;
  wire       [2:0]    _zz_59;
  wire       [1:0]    _zz_LsuL1Plugin_logic_shared_write_payload_data_dirty;
  wire       [0:0]    _zz_when;
  wire       [0:0]    _zz_LsuL1Plugin_logic_waysWrite_tag_fault;
  reg        [19:0]   _zz__zz_LsuL1Plugin_logic_waysWrite_tag_address;
  reg                 _zz_LsuL1Plugin_logic_waysWrite_tag_fault_1;
  reg        [19:0]   _zz_LsuL1Plugin_logic_writeback_push_payload_address;
  wire       [0:0]    _zz_LsuL1Plugin_logic_shared_write_payload_data_plru_0_1;
  wire       [64:0]   _zz_execute_ctrl2_down_MUL_SRC1_lane0;
  wire       [64:0]   _zz_execute_ctrl2_down_MUL_SRC2_lane0;
  wire       [76:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_6_lane0;
  wire       [31:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_6_lane0_1;
  wire       [17:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_6_lane0_2;
  wire       [13:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_6_lane0_3;
  wire       [76:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_7_lane0;
  wire       [31:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_7_lane0_1;
  wire       [13:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_7_lane0_2;
  wire       [17:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_7_lane0_3;
  wire       [59:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_10_lane0;
  wire       [31:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_10_lane0_1;
  wire       [17:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_10_lane0_2;
  wire       [13:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_10_lane0_3;
  wire       [59:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_11_lane0;
  wire       [31:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_11_lane0_1;
  wire       [13:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_11_lane0_2;
  wire       [17:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_11_lane0_3;
  wire       [42:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_13_lane0;
  wire       [31:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_13_lane0_1;
  wire       [17:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_13_lane0_2;
  wire       [13:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_13_lane0_3;
  wire       [42:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_14_lane0;
  wire       [31:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_14_lane0_1;
  wire       [13:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_14_lane0_2;
  wire       [17:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_14_lane0_3;
  wire       [25:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_15_lane0;
  wire       [27:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_15_lane0_1;
  wire       [13:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_15_lane0_2;
  wire       [13:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_15_lane0_3;
  wire       [63:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_7;
  wire       [63:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_8;
  wire       [63:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_9;
  wire       [63:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_10;
  wire       [63:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_11;
  wire       [63:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_12;
  wire       [63:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_13;
  wire       [63:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_14;
  wire       [63:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_15;
  wire       [63:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_16;
  wire       [63:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_17;
  wire       [63:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_18;
  wire       [46:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_7;
  wire       [46:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_8;
  wire       [46:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_9;
  wire       [46:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_10;
  wire       [46:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_11;
  wire       [46:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_12;
  wire       [46:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_13;
  wire       [46:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_14;
  wire       [46:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_15;
  wire       [46:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_16;
  wire       [46:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_17;
  wire       [46:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_18;
  wire       [25:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_7;
  wire       [25:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_8;
  wire       [25:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_9;
  wire       [25:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_10;
  wire       [25:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_11;
  wire       [25:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_12;
  wire       [25:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_13;
  wire       [25:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_14;
  wire       [25:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_15;
  wire       [25:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_16;
  wire       [25:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_17;
  wire       [25:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_18;
  wire       [63:0]   _zz_execute_ctrl2_down_RsUnsignedPlugin_RS1_UNSIGNED_lane0;
  wire       [0:0]    _zz_execute_ctrl2_down_RsUnsignedPlugin_RS1_UNSIGNED_lane0_1;
  wire       [63:0]   _zz_execute_ctrl2_down_RsUnsignedPlugin_RS2_UNSIGNED_lane0;
  wire       [0:0]    _zz_execute_ctrl2_down_RsUnsignedPlugin_RS2_UNSIGNED_lane0_1;
  wire       [63:0]   _zz_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0_1;
  wire       [63:0]   _zz_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0_2;
  wire       [0:0]    _zz_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0_3;
  wire       [21:0]   _zz_FetchL1Plugin_logic_ways_0_mem_port;
  wire                _zz_FetchL1Plugin_logic_ways_0_mem_port_1;
  wire       [21:0]   _zz_FetchL1Plugin_logic_ways_1_mem_port;
  wire                _zz_FetchL1Plugin_logic_ways_1_mem_port_1;
  wire                _zz_when_1;
  reg        [31:0]   _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_0;
  wire       [0:0]    _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_0_1;
  reg        [31:0]   _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_1;
  wire       [0:0]    _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_1_1;
  wire       [26:0]   _zz_FetchL1Plugin_logic_hits_w_0_indirect_bypassHits;
  wire       [26:0]   _zz_FetchL1Plugin_logic_hits_w_0_indirect_bypassHits_1;
  wire       [26:0]   _zz_FetchL1Plugin_logic_hits_w_1_indirect_bypassHits;
  wire       [26:0]   _zz_FetchL1Plugin_logic_hits_w_1_indirect_bypassHits_1;
  wire       [0:0]    _zz_FetchL1Plugin_logic_ctrl_dataAccessFault;
  wire       [0:0]    _zz_FetchL1Plugin_logic_plru_write_payload_data_0;
  wire       [3:0]    _zz_GSharePlugin_logic_mem_banks_0_port;
  wire                _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_1;
  wire       [0:0]    _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_2;
  wire       [4:0]    _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_3;
  wire       [12:0]   _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_4;
  wire       [11:0]   _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_5;
  wire       [1:0]    _zz_BtbPlugin_logic_ras_ptr_push;
  wire       [1:0]    _zz_BtbPlugin_logic_ras_ptr_push_1;
  wire       [0:0]    _zz_BtbPlugin_logic_ras_ptr_push_2;
  wire       [1:0]    _zz_BtbPlugin_logic_ras_ptr_push_3;
  wire       [0:0]    _zz_BtbPlugin_logic_ras_ptr_push_4;
  wire       [1:0]    _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue;
  wire       [1:0]    _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_1;
  wire       [0:0]    _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_2;
  wire       [1:0]    _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_3;
  wire       [0:0]    _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_4;
  wire       [37:0]   _zz_BtbPlugin_logic_ras_mem_stack_port;
  wire       [57:0]   _zz_BtbPlugin_logic_mem_port;
  wire       [63:0]   _zz_WhiteboxerPlugin_logic_decodes_0_pc;
  wire       [38:0]   _zz_WhiteboxerPlugin_logic_decodes_0_pc_1;
  wire       [0:0]    _zz_FetchL1Plugin_pmaBuilder_onTransfers_0_addressHit;
  wire       [0:0]    _zz_FetchL1Plugin_logic_ctrl_pmaPort_rsp_io_1;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_commitCount;
  wire       [0:0]    _zz_PerformanceCounterPlugin_logic_commitCount_1;
  wire       [0:0]    _zz_PerformanceCounterPlugin_logic_eventInstructions_0;
  wire       [7:0]    _zz_PerformanceCounterPlugin_logic_counters_cycle_value;
  wire       [0:0]    _zz_PerformanceCounterPlugin_logic_counters_cycle_value_1;
  wire       [7:0]    _zz_PerformanceCounterPlugin_logic_counters_instret_value_1;
  wire       [63:0]   _zz_LsuPlugin_logic_onAddress0_ls_port_payload_address;
  wire       [11:0]   _zz_LsuPlugin_logic_onAddress0_ls_storeId;
  wire       [0:0]    _zz_LsuPlugin_logic_onAddress0_ls_storeId_1;
  wire       [12:0]   _zz_LsuPlugin_logic_onAddress0_flush_port_payload_address;
  wire       [63:0]   _zz_LsuPlugin_logic_onPma_addressExtension;
  wire       [24:0]   _zz__zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0;
  wire                _zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0_1;
  wire                _zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0_2;
  wire       [0:0]    _zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0_3;
  wire       [18:0]   _zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0_4;
  wire                _zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0_5;
  wire                _zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0_6;
  wire       [0:0]    _zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0_7;
  wire       [10:0]   _zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0_8;
  wire                _zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0_9;
  wire                _zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0_10;
  wire       [0:0]    _zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0_11;
  wire       [2:0]    _zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0_12;
  reg        [7:0]    _zz_LsuPlugin_logic_onCtrl_loadData_shifted;
  wire       [2:0]    _zz_LsuPlugin_logic_onCtrl_loadData_shifted_1;
  reg        [7:0]    _zz_LsuPlugin_logic_onCtrl_loadData_shifted_2;
  wire       [1:0]    _zz_LsuPlugin_logic_onCtrl_loadData_shifted_3;
  reg        [7:0]    _zz_LsuPlugin_logic_onCtrl_loadData_shifted_4;
  wire       [0:0]    _zz_LsuPlugin_logic_onCtrl_loadData_shifted_5;
  reg        [7:0]    _zz_LsuPlugin_logic_onCtrl_loadData_shifted_6;
  wire       [0:0]    _zz_LsuPlugin_logic_onCtrl_loadData_shifted_7;
  wire       [63:0]   _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub;
  wire       [63:0]   _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_1;
  wire       [63:0]   _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_2;
  wire       [63:0]   _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_3;
  wire       [63:0]   _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_4;
  wire       [1:0]    _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_5;
  wire       [2:0]    _zz_LsuPlugin_logic_trapPort_payload_code;
  wire                _zz_execute_ctrl4_down_LsuL1_ABORD_lane0;
  wire       [5:0]    _zz_LsuPlugin_logic_flusher_cmdCounter;
  wire       [31:0]   _zz__zz_execute_ctrl1_down_early0_SrcPlugin_SRC1_lane0;
  wire       [11:0]   _zz__zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0;
  wire       [38:0]   _zz__zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0_1;
  wire       [11:0]   _zz__zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0_2;
  wire       [63:0]   _zz_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0;
  wire       [63:0]   _zz_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0_1;
  wire       [63:0]   _zz_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0_2;
  wire       [0:0]    _zz_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0_3;
  wire       [20:0]   _zz_early0_BranchPlugin_pcCalc_target_b;
  wire       [11:0]   _zz_early0_BranchPlugin_pcCalc_target_b_1;
  wire       [12:0]   _zz_early0_BranchPlugin_pcCalc_target_b_2;
  wire       [63:0]   _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0;
  wire       [63:0]   _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0_1;
  wire       [63:0]   _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0_2;
  wire       [38:0]   _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0;
  wire       [2:0]    _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0_1;
  wire       [38:0]   _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0;
  wire       [1:0]    _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0_1;
  reg        [1:0]    _zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK;
  wire       [0:0]    _zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK_1;
  reg        [1:0]    _zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK_2;
  wire       [1:0]    _zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_LAST;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_redo_4;
  wire       [4:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_19;
  wire       [0:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_20;
  wire                _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_21;
  wire       [31:0]   _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_22;
  wire       [11:0]   _zz__zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_18;
  wire       [5:0]    _zz__zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_18_1;
  reg        [31:0]   _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_23;
  wire       [1:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_24;
  reg        [2:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_25;
  wire       [2:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_26;
  wire       [6:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_27;
  wire       [4:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_28;
  wire                _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_29;
  wire       [4:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_30;
  wire       [11:0]   _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_31;
  wire       [11:0]   _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_32;
  wire       [11:0]   _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_33;
  wire       [11:0]   _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_34;
  wire       [1:0]    _zz__zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_5;
  wire       [38:0]   _zz_early0_EnvPlugin_logic_trapPort_payload_tval;
  wire       [31:0]   _zz_early0_EnvPlugin_logic_trapPort_payload_tval_1;
  wire       [3:0]    _zz_early0_EnvPlugin_logic_trapPort_payload_code;
  wire       [31:0]   _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_napot_MATCH;
  wire       [19:0]   _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_tor_BIGGER;
  wire       [31:0]   _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_napot_MATCH;
  wire       [19:0]   _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_tor_BIGGER;
  wire       [31:0]   _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_napot_MATCH;
  wire       [19:0]   _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_tor_BIGGER;
  wire       [31:0]   _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_napot_MATCH;
  wire       [19:0]   _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_tor_BIGGER;
  wire       [0:0]    _zz_fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_ACCESS_FAULT_4;
  wire       [0:0]    _zz_fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_ACCESS_FAULT_5;
  wire       [31:0]   _zz_execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_0_napot_MATCH_lane0;
  wire       [19:0]   _zz_execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_0_tor_BIGGER_lane0;
  wire       [31:0]   _zz_execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_1_napot_MATCH_lane0;
  wire       [19:0]   _zz_execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_1_tor_BIGGER_lane0;
  wire       [31:0]   _zz_execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_2_napot_MATCH_lane0;
  wire       [19:0]   _zz_execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_2_tor_BIGGER_lane0;
  wire       [31:0]   _zz_execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_3_napot_MATCH_lane0;
  wire       [19:0]   _zz_execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_3_tor_BIGGER_lane0;
  wire       [0:0]    _zz_execute_ctrl4_down_LsuPlugin_logic_pmpPort_ACCESS_FAULT_lane0_4;
  wire       [0:0]    _zz_execute_ctrl4_down_LsuPlugin_logic_pmpPort_ACCESS_FAULT_lane0_5;
  wire       [0:0]    _zz_LsuPlugin_pmaBuilder_l1_onTransfers_0_addressHit;
  wire       [0:0]    _zz_LsuPlugin_logic_onPma_cached_rsp_io_1;
  wire       [0:0]    _zz_LsuPlugin_pmaBuilder_io_onTransfers_0_addressHit;
  wire       [31:0]   _zz_LsuPlugin_logic_onPma_io_rsp_fault;
  wire       [31:0]   _zz_LsuPlugin_logic_onPma_io_rsp_fault_1;
  wire       [31:0]   _zz_LsuPlugin_logic_onPma_io_rsp_fault_2;
  wire                _zz_LsuPlugin_logic_onPma_io_rsp_fault_3;
  wire       [0:0]    _zz_LsuPlugin_logic_onPma_io_rsp_fault_4;
  wire       [3:0]    _zz_LsuPlugin_logic_onPma_io_rsp_fault_5;
  wire       [0:0]    _zz_LsuPlugin_logic_onPma_io_rsp_io;
  wire       [63:0]   _zz_early0_BranchPlugin_logic_alu_expectedMsb;
  wire       [24:0]   _zz__zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0;
  wire                _zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0_1;
  wire                _zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0_2;
  wire       [0:0]    _zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0_3;
  wire       [18:0]   _zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0_4;
  wire                _zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0_5;
  wire                _zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0_6;
  wire       [0:0]    _zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0_7;
  wire       [10:0]   _zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0_8;
  wire                _zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0_9;
  wire                _zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0_10;
  wire       [0:0]    _zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0_11;
  wire       [2:0]    _zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0_12;
  wire       [12:0]   _zz_early0_BranchPlugin_logic_jumpLogic_history_shifter_1;
  wire       [12:0]   _zz_early0_BranchPlugin_logic_jumpLogic_history_shifter_2;
  wire       [63:0]   _zz_early0_BranchPlugin_logic_wb_payload;
  wire       [38:0]   _zz_early0_BranchPlugin_logic_wb_payload_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_RS1_ENABLE_0;
  wire       [31:0]   _zz_decode_ctrls_1_down_RS1_ENABLE_0_1;
  wire       [31:0]   _zz_decode_ctrls_1_down_RS1_ENABLE_0_2;
  wire       [4:0]    _zz_decode_ctrls_1_down_RS1_PHYS_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_RS2_ENABLE_0;
  wire       [4:0]    _zz_decode_ctrls_1_down_RS2_PHYS_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_RD_ENABLE_0;
  wire       [31:0]   _zz_decode_ctrls_1_down_RD_ENABLE_0_1;
  wire       [31:0]   _zz_decode_ctrls_1_down_RD_ENABLE_0_2;
  wire       [31:0]   _zz_decode_ctrls_1_down_RD_ENABLE_0_3;
  wire       [31:0]   _zz_decode_ctrls_1_down_RD_ENABLE_0_4;
  wire       [31:0]   _zz_decode_ctrls_1_down_RD_ENABLE_0_5;
  wire       [4:0]    _zz_decode_ctrls_1_down_RD_PHYS_0;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_1;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_2;
  wire                _zz_decode_ctrls_1_down_Decode_LEGAL_0_3;
  wire       [0:0]    _zz_decode_ctrls_1_down_Decode_LEGAL_0_4;
  wire       [22:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_5;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_6;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_7;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_8;
  wire                _zz_decode_ctrls_1_down_Decode_LEGAL_0_9;
  wire       [0:0]    _zz_decode_ctrls_1_down_Decode_LEGAL_0_10;
  wire       [16:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_11;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_12;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_13;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_14;
  wire                _zz_decode_ctrls_1_down_Decode_LEGAL_0_15;
  wire       [0:0]    _zz_decode_ctrls_1_down_Decode_LEGAL_0_16;
  wire       [10:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_17;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_18;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_19;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_20;
  wire                _zz_decode_ctrls_1_down_Decode_LEGAL_0_21;
  wire       [0:0]    _zz_decode_ctrls_1_down_Decode_LEGAL_0_22;
  wire       [4:0]    _zz_decode_ctrls_1_down_Decode_LEGAL_0_23;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_24;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_25;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_26;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_27;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_28;
  wire       [0:0]    _zz_DecoderPlugin_logic_laneLogic_0_fixer_isJb;
  wire       [38:0]   _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice;
  wire       [1:0]    _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice_1;
  wire       [1:0]    _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice_2;
  wire       [11:0]   _zz_CsrRamPlugin_csrMapper_ramAddress_1;
  wire       [11:0]   _zz_CsrRamPlugin_csrMapper_ramAddress_2;
  wire       [11:0]   _zz_CsrRamPlugin_csrMapper_ramAddress_3;
  wire       [11:0]   _zz_CsrRamPlugin_csrMapper_ramAddress_4;
  wire                _zz_CsrRamPlugin_csrMapper_ramAddress_5;
  wire       [0:0]    _zz_CsrRamPlugin_csrMapper_ramAddress_6;
  wire       [11:0]   _zz_CsrRamPlugin_csrMapper_ramAddress_7;
  wire       [0:0]    _zz_CsrRamPlugin_csrMapper_ramAddress_8;
  wire       [11:0]   _zz_CsrRamPlugin_csrMapper_ramAddress_9;
  wire                _zz_CsrRamPlugin_csrMapper_ramAddress_10;
  wire       [0:0]    _zz_CsrRamPlugin_csrMapper_ramAddress_11;
  wire       [11:0]   _zz_CsrRamPlugin_csrMapper_ramAddress_12;
  wire       [0:0]    _zz_CsrRamPlugin_csrMapper_ramAddress_13;
  wire       [11:0]   _zz_CsrRamPlugin_csrMapper_ramAddress_14;
  wire                _zz_GSharePlugin_logic_onLearn_hash_1;
  wire       [0:0]    _zz_GSharePlugin_logic_onLearn_hash_2;
  wire       [4:0]    _zz_GSharePlugin_logic_onLearn_hash_3;
  wire       [12:0]   _zz_GSharePlugin_logic_onLearn_hash_4;
  wire       [11:0]   _zz_GSharePlugin_logic_onLearn_hash_5;
  wire       [36:0]   _zz_BtbPlugin_logic_memWrite_payload_address;
  wire       [0:0]    _zz_decode_ctrls_1_down_AguPlugin_CLEAN_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_AguPlugin_CLEAN_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_AguPlugin_INVALIDATE_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_AguPlugin_INVALIDATE_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_2;
  wire       [0:0]    _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_3;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0_2;
  wire       [36:0]   _zz_BtbPlugin_logic_memWrite_payload_address_1;
  wire       [36:0]   _zz_BtbPlugin_logic_memRead_cmd_payload;
  wire       [38:0]   _zz_BtbPlugin_logic_ras_write_payload_data;
  wire       [39:0]   _zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception;
  wire       [39:0]   _zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception_1;
  wire       [39:0]   _zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception_2;
  wire       [39:0]   _zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception_3;
  wire       [1:0]    _zz_TrapPlugin_logic_harts_0_trap_pending_slices;
  wire       [38:0]   _zz_TrapPlugin_logic_harts_0_trap_fsm_jumpTarget;
  wire       [2:0]    _zz_TrapPlugin_logic_harts_0_trap_fsm_jumpTarget_1;
  wire       [38:0]   _zz_PcPlugin_logic_harts_0_self_pc;
  wire       [2:0]    _zz_PcPlugin_logic_harts_0_self_pc_1;
  wire       [0:0]    _zz_PcPlugin_logic_harts_0_aggregator_fault;
  wire       [0:0]    _zz_PcPlugin_logic_harts_0_aggregator_fault_1_1;
  wire       [46:0]   _zz_FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_0_port;
  wire                _zz_FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_0_port_1;
  wire       [46:0]   _zz_FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_1_port;
  wire                _zz_FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_1_port_1;
  wire       [28:0]   _zz_FetchL1Plugin_logic_translationStorage_logic_sl_1_ways_0_port;
  wire                _zz_FetchL1Plugin_logic_translationStorage_logic_sl_1_ways_0_port_1;
  wire       [46:0]   _zz_LsuPlugin_logic_translationStorage_logic_sl_0_ways_0_port;
  wire                _zz_LsuPlugin_logic_translationStorage_logic_sl_0_ways_0_port_1;
  wire       [46:0]   _zz_LsuPlugin_logic_translationStorage_logic_sl_0_ways_1_port;
  wire                _zz_LsuPlugin_logic_translationStorage_logic_sl_0_ways_1_port_1;
  wire       [46:0]   _zz_LsuPlugin_logic_translationStorage_logic_sl_0_ways_2_port;
  wire                _zz_LsuPlugin_logic_translationStorage_logic_sl_0_ways_2_port_1;
  wire       [1:0]    _zz_LsuPlugin_logic_translationStorage_logic_sl_0_allocId_valueNext;
  wire       [0:0]    _zz_LsuPlugin_logic_translationStorage_logic_sl_0_allocId_valueNext_1;
  wire       [28:0]   _zz_LsuPlugin_logic_translationStorage_logic_sl_1_ways_0_port;
  wire                _zz_LsuPlugin_logic_translationStorage_logic_sl_1_ways_0_port_1;
  wire       [0:0]    _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_4;
  wire       [0:0]    _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowRead;
  wire       [0:0]    _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowWrite;
  wire       [0:0]    _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowUser;
  wire       [19:0]   _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated;
  wire       [11:0]   _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_1;
  wire       [19:0]   _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_2;
  wire       [11:0]   _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_3;
  wire       [19:0]   _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_4;
  wire       [11:0]   _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_5;
  wire       [10:0]   _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_6;
  wire       [20:0]   _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_7;
  wire       [0:0]    _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_3;
  wire       [0:0]    _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowRead;
  wire       [0:0]    _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowWrite;
  wire       [0:0]    _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowUser;
  wire       [11:0]   _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineTranslated;
  wire       [11:0]   _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineTranslated_1;
  wire       [25:0]   _zz_MmuPlugin_logic_refill_load_nextLevelBase;
  wire       [53:0]   _zz_bits_pte_ppn;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_0_1;
  wire       [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_0_2;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_1_1;
  wire       [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_1_2;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_2_1;
  wire       [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_2_2;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_3_1;
  wire       [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_3_2;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_4_1;
  wire       [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_4_2;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_5_1;
  wire       [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_5_2;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_6_1;
  wire       [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_6_2;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_7_1;
  wire       [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_7_2;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_8_1;
  wire       [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_8_2;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_9_1;
  wire       [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_9_2;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_10_1;
  wire       [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_10_2;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_11_1;
  wire       [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_11_2;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_12_1;
  wire       [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_12_2;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_13_1;
  wire       [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_13_2;
  wire       [6:0]    _zz_PerformanceCounterPlugin_logic_fsm_calc_a;
  wire       [64:0]   _zz_PerformanceCounterPlugin_logic_fsm_calc_sum;
  wire       [8:0]    _zz_PerformanceCounterPlugin_logic_fsm_calc_sum_1;
  wire       [1:0]    _zz_PerformanceCounterPlugin_logic_flusher_hits_ohFirst_masked;
  wire                _zz_fetch_logic_flushes_0_doIt;
  wire                _zz_fetch_logic_flushes_0_doIt_1;
  wire                _zz_fetch_logic_flushes_0_doIt_2;
  wire       [11:0]   _zz_COMB_CSR_PmpPlugin_logic_allFilter;
  wire                _zz_COMB_CSR_PmpPlugin_logic_allFilter_1;
  wire       [0:0]    _zz_COMB_CSR_PmpPlugin_logic_allFilter_2;
  wire       [10:0]   _zz_COMB_CSR_PmpPlugin_logic_allFilter_3;
  wire       [11:0]   _zz_COMB_CSR_PmpPlugin_logic_allFilter_4;
  wire                _zz_COMB_CSR_PmpPlugin_logic_allFilter_5;
  wire       [0:0]    _zz_COMB_CSR_PmpPlugin_logic_allFilter_6;
  wire       [2:0]    _zz_COMB_CSR_PmpPlugin_logic_allFilter_7;
  wire       [11:0]   _zz_COMB_CSR_UNAMED_1;
  wire                _zz_COMB_CSR_UNAMED_1_1;
  wire       [0:0]    _zz_COMB_CSR_UNAMED_1_2;
  wire       [77:0]   _zz_COMB_CSR_UNAMED_1_3;
  wire       [11:0]   _zz_COMB_CSR_UNAMED_1_4;
  wire                _zz_COMB_CSR_UNAMED_1_5;
  wire       [0:0]    _zz_COMB_CSR_UNAMED_1_6;
  wire       [69:0]   _zz_COMB_CSR_UNAMED_1_7;
  wire       [11:0]   _zz_COMB_CSR_UNAMED_1_8;
  wire                _zz_COMB_CSR_UNAMED_1_9;
  wire       [0:0]    _zz_COMB_CSR_UNAMED_1_10;
  wire       [61:0]   _zz_COMB_CSR_UNAMED_1_11;
  wire       [11:0]   _zz_COMB_CSR_UNAMED_1_12;
  wire                _zz_COMB_CSR_UNAMED_1_13;
  wire       [0:0]    _zz_COMB_CSR_UNAMED_1_14;
  wire       [53:0]   _zz_COMB_CSR_UNAMED_1_15;
  wire       [11:0]   _zz_COMB_CSR_UNAMED_1_16;
  wire                _zz_COMB_CSR_UNAMED_1_17;
  wire       [0:0]    _zz_COMB_CSR_UNAMED_1_18;
  wire       [45:0]   _zz_COMB_CSR_UNAMED_1_19;
  wire       [11:0]   _zz_COMB_CSR_UNAMED_1_20;
  wire                _zz_COMB_CSR_UNAMED_1_21;
  wire       [0:0]    _zz_COMB_CSR_UNAMED_1_22;
  wire       [37:0]   _zz_COMB_CSR_UNAMED_1_23;
  wire       [11:0]   _zz_COMB_CSR_UNAMED_1_24;
  wire                _zz_COMB_CSR_UNAMED_1_25;
  wire       [0:0]    _zz_COMB_CSR_UNAMED_1_26;
  wire       [29:0]   _zz_COMB_CSR_UNAMED_1_27;
  wire       [11:0]   _zz_COMB_CSR_UNAMED_1_28;
  wire                _zz_COMB_CSR_UNAMED_1_29;
  wire       [0:0]    _zz_COMB_CSR_UNAMED_1_30;
  wire       [21:0]   _zz_COMB_CSR_UNAMED_1_31;
  wire       [11:0]   _zz_COMB_CSR_UNAMED_1_32;
  wire                _zz_COMB_CSR_UNAMED_1_33;
  wire       [0:0]    _zz_COMB_CSR_UNAMED_1_34;
  wire       [13:0]   _zz_COMB_CSR_UNAMED_1_35;
  wire       [11:0]   _zz_COMB_CSR_UNAMED_1_36;
  wire                _zz_COMB_CSR_UNAMED_1_37;
  wire       [0:0]    _zz_COMB_CSR_UNAMED_1_38;
  wire       [5:0]    _zz_COMB_CSR_UNAMED_1_39;
  wire       [11:0]   _zz_COMB_CSR_CsrRamPlugin_csrMapper_selFilter;
  wire                _zz_COMB_CSR_CsrRamPlugin_csrMapper_selFilter_1;
  wire       [0:0]    _zz_COMB_CSR_CsrRamPlugin_csrMapper_selFilter_2;
  wire       [2:0]    _zz_COMB_CSR_CsrRamPlugin_csrMapper_selFilter_3;
  wire       [0:0]    _zz_CsrAccessPlugin_logic_fsm_inject_implemented;
  wire       [28:0]   _zz_CsrAccessPlugin_logic_fsm_inject_implemented_1;
  wire       [0:0]    _zz_CsrAccessPlugin_logic_fsm_inject_implemented_2;
  wire       [17:0]   _zz_CsrAccessPlugin_logic_fsm_inject_implemented_3;
  wire       [0:0]    _zz_CsrAccessPlugin_logic_fsm_inject_implemented_4;
  wire       [6:0]    _zz_CsrAccessPlugin_logic_fsm_inject_implemented_5;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_32;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_33;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_34;
  wire       [19:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_35;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_36;
  wire       [18:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_37;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_38;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_39;
  wire       [19:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_40;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_41;
  wire       [18:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_42;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_43;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_44;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_45;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_46;
  wire       [43:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_47;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_48;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_49;
  wire       [43:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_50;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_51;
  wire       [29:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_52;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_53;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_54;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_55;
  wire       [9:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_56;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_57;
  wire       [0:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_58;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_59;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_60;
  wire       [1:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_61;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_62;
  wire       [2:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_63;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_64;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_65;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_66;
  wire       [4:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_67;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_68;
  wire       [7:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_69;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_70;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_71;
  wire       [29:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_72;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_73;
  wire       [9:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_74;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_75;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_76;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_77;
  wire       [8:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_78;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_79;
  wire       [9:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_80;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_81;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_82;
  wire       [10:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_83;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_84;
  wire       [12:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_85;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_86;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_87;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_88;
  wire       [15:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_89;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_90;
  wire       [29:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_91;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_92;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_93;
  wire       [9:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_94;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_95;
  wire       [16:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_96;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_97;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_98;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_99;
  wire       [17:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_100;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_101;
  wire       [18:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_102;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_103;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_104;
  wire       [20:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_105;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_106;
  wire       [23:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_107;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_108;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_109;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_110;
  wire       [29:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_111;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_112;
  wire       [9:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_113;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_114;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_115;
  wire       [24:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_116;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_117;
  wire       [25:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_118;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_119;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_120;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_121;
  wire       [26:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_122;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_123;
  wire       [28:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_124;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_125;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_126;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_127;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_128;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_129;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_130;
  wire       [5:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_131;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_132;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_133;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_134;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_135;
  wire       [7:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_136;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_137;
  wire       [3:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_138;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_139;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_140;
  wire       [12:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_141;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_142;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_143;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_144;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_145;
  wire       [17:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_146;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_147;
  wire       [14:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_148;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_149;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_150;
  wire       [33:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_151;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_152;
  wire       [35:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_153;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_154;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_155;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_156;
  wire       [22:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_157;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_158;
  wire       [20:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_159;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_160;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_161;
  wire       [21:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_162;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_163;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_164;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_165;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_166;
  wire       [3:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_167;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_168;
  wire       [11:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_169;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_170;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_171;
  wire       [7:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_172;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_173;
  wire       [3:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_174;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_175;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_176;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_177;
  wire       [11:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_178;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_179;
  wire       [7:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_180;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_181;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_182;
  wire       [3:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_183;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_184;
  wire       [0:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_185;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_186;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_187;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_188;
  wire       [3:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_189;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_190;
  wire       [8:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_191;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_192;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_193;
  wire       [9:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_194;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_195;
  wire       [12:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_196;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_197;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_198;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_199;
  wire       [13:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_200;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_201;
  wire       [15:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_202;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_203;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_204;
  wire       [9:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_205;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_206;
  wire       [5:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_207;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_208;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_209;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_210;
  wire       [1:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_211;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_212;
  wire       [0:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_213;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_214;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_215;
  wire       [19:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_216;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_217;
  wire       [1:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_218;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_219;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_220;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_221;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_222;
  wire       [3:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_223;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_224;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_225;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_226;
  wire       [8:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_227;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_228;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_229;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_230;
  wire       [5:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_231;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_232;
  wire       [1:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_233;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_234;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_235;
  wire       [8:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_236;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_237;
  wire       [5:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_238;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_239;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_240;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_241;
  wire       [1:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_242;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_243;
  wire       [33:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_244;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_245;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_246;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_247;
  wire       [14:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_248;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_249;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_250;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_251;
  wire       [9:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_252;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_253;
  wire       [5:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_254;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_255;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_256;
  wire       [1:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_257;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_258;
  wire       [9:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_259;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_260;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_261;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_262;
  wire       [1:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_263;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_264;
  wire       [9:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_265;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_266;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_267;
  wire       [5:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_268;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_269;
  wire       [1:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_270;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_271;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_272;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_273;
  wire       [9:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_274;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_275;
  wire       [5:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_276;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_277;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_278;
  wire       [5:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_279;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_280;
  wire       [1:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_281;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_282;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_283;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_284;
  wire       [0:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_285;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_286;
  wire       [19:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_287;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_288;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_289;
  wire       [0:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_290;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_291;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_292;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_293;
  wire       [0:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_294;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_295;
  wire       [0:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_296;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_297;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_298;
  wire       [2:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_299;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_300;
  wire       [2:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_301;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_302;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_303;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_304;
  wire       [2:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_305;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_306;
  wire       [5:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_307;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_308;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_309;
  wire       [6:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_310;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_311;
  wire       [5:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_312;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_313;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_314;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_315;
  wire       [6:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_316;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_317;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_318;
  wire       [13:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_319;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_320;
  wire       [13:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_321;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_322;
  wire       [13:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_323;
  wire       [63:0]   _zz_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask;
  wire       [4:0]    _zz_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask_1;
  wire       [3:0]    _zz_CsrRamPlugin_logic_writeLogic_hits_ohFirst_masked;
  wire       [2:0]    _zz_CsrRamPlugin_logic_readLogic_hits_ohFirst_masked;
  reg        [3:0]    _zz_CsrRamPlugin_logic_readLogic_port_cmd_payload;
  wire       [4:0]    _zz_CsrRamPlugin_logic_flush_counter;
  wire       [0:0]    _zz_CsrRamPlugin_logic_flush_counter_1;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0_2;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_BarrelShifterPlugin_SEL_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_BarrelShifterPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_BranchPlugin_SEL_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_BranchPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_MulPlugin_SEL_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_MulPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_DivPlugin_SEL_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_DivPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_EnvPlugin_SEL_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_EnvPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_MulPlugin_HIGH_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_MulPlugin_HIGH_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_CsrAccessPlugin_SEL_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_CsrAccessPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_AguPlugin_SEL_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_AguPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_LsuPlugin_logic_FENCE_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_LsuPlugin_logic_FENCE_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_COMPLETION_AT_2_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_COMPLETION_AT_2_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_COMPLETION_AT_4_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_COMPLETION_AT_4_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_COMPLETION_AT_3_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_COMPLETION_AT_3_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_4;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_5;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_4;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_5;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0_3;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0_4;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0_2;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_SLTX_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_SLTX_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_SrcStageables_REVERT_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_SrcStageables_REVERT_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_SrcStageables_ZERO_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_SrcStageables_ZERO_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_SIGNED_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_SIGNED_lane0_1;
  wire       [31:0]   _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
  wire       [31:0]   _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0_1;
  wire       [31:0]   _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0_2;
  wire                _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0_3;
  wire       [31:0]   _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0_4;
  wire       [31:0]   _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0_5;
  wire       [31:0]   _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0_6;
  wire                _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0_7;
  wire                _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0_8;
  wire       [0:0]    _zz_execute_ctrl1_down_BYPASSED_AT_2_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_BYPASSED_AT_2_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_BYPASSED_AT_3_lane0_3;
  wire       [0:0]    _zz_execute_ctrl1_down_BYPASSED_AT_3_lane0_4;
  wire       [0:0]    _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_SrcStageables_UNSIGNED_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_SrcStageables_UNSIGNED_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0_2;
  wire       [0:0]    _zz_execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_BarrelShifterPlugin_IS_W_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_BarrelShifterPlugin_IS_W_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_BarrelShifterPlugin_IS_W_RIGHT_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_BarrelShifterPlugin_IS_W_RIGHT_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_RsUnsignedPlugin_RS1_SIGNED_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_RsUnsignedPlugin_RS1_SIGNED_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0_2;
  wire       [0:0]    _zz_execute_ctrl1_down_DivPlugin_REM_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_DivPlugin_REM_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_RsUnsignedPlugin_IS_W_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_RsUnsignedPlugin_IS_W_lane0_2;
  wire       [0:0]    _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_IMM_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_IMM_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0_2;
  wire       [0:0]    _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0_2;
  wire       [0:0]    _zz_execute_ctrl1_down_AguPlugin_LOAD_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_AguPlugin_LOAD_lane0_2;
  wire       [0:0]    _zz_execute_ctrl1_down_AguPlugin_STORE_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_AguPlugin_STORE_lane0_2;
  wire       [0:0]    _zz_execute_ctrl1_down_AguPlugin_ATOMIC_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_AguPlugin_ATOMIC_lane0_2;
  wire       [0:0]    _zz_execute_ctrl1_down_AguPlugin_FLOAT_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_AguPlugin_FLOAT_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_AguPlugin_CLEAN_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_AguPlugin_CLEAN_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_AguPlugin_INVALIDATE_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_AguPlugin_INVALIDATE_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_LsuPlugin_logic_LSU_PREFETCH_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_LsuPlugin_logic_LSU_PREFETCH_lane0_1;
  wire       [31:0]   _zz__zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2;
  wire       [31:0]   _zz__zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_1;
  wire       [31:0]   _zz__zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_2;
  wire       [31:0]   _zz__zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_3;
  wire                _zz__zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_4;
  wire                _zz__zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_5;
  wire                _zz_when_ExecuteLanePlugin_l306_2;
  wire                _zz_when_ExecuteLanePlugin_l306_2_1;
  wire                _zz_when_ExecuteLanePlugin_l306_2_2;
  wire                _zz_when_ExecuteLanePlugin_l306_2_3;
  wire       [31:0]   _zz_WhiteboxerPlugin_logic_csr_access_payload_address;
  reg        [0:0]    _zz_WhiteboxerPlugin_logic_perf_candidatesCount;
  wire       [0:0]    _zz_WhiteboxerPlugin_logic_perf_candidatesCount_1;
  reg        [0:0]    _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCount;
  wire       [0:0]    _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCount_1;
  wire       [59:0]   _zz__zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_1;
  wire       [0:0]    _zz__zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_1_1;
  wire       [59:0]   _zz__zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_1;
  wire       [0:0]    _zz__zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_1_1;
  wire       [59:0]   _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_1;
  wire       [0:0]    _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_1_1;
  wire       [59:0]   _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_1;
  wire       [0:0]    _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_1_1;
  wire       [59:0]   _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_1;
  wire       [0:0]    _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_1_1;
  wire       [59:0]   _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_1;
  wire       [0:0]    _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_1_1;
  wire       [63:0]   _zz_TrapPlugin_logic_harts_0_crsPorts_write_data;
  wire       [38:0]   _zz_TrapPlugin_logic_harts_0_crsPorts_write_data_1;
  wire       [63:0]   _zz_TrapPlugin_logic_harts_0_crsPorts_write_data_2;
  wire       [38:0]   _zz_TrapPlugin_logic_harts_0_crsPorts_write_data_3;
  wire       [63:0]   _zz_TrapPlugin_logic_harts_0_crsPorts_write_data_4;
  wire       [38:0]   _zz_TrapPlugin_logic_harts_0_crsPorts_write_data_5;
  wire       [63:0]   _zz_TrapPlugin_logic_harts_0_trap_pcPort_payload_pc;
  wire       [63:0]   _zz_TrapPlugin_logic_harts_0_trap_pcPort_payload_pc_1;
  wire       [55:0]   _zz_MmuPlugin_logic_refill_load_address;
  wire       [1:0]    _zz_FetchL1Plugin_logic_translationStorage_logic_sl_0_write_mask;
  wire       [43:0]   _zz_FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_physicalAddress;
  wire       [3:0]    _zz_LsuPlugin_logic_translationStorage_logic_sl_0_write_mask;
  wire       [3:0]    _zz_LsuPlugin_logic_translationStorage_logic_sl_0_write_mask_1;
  wire       [43:0]   _zz_LsuPlugin_logic_translationStorage_logic_sl_0_write_data_physicalAddress;
  wire       [34:0]   _zz_FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_physicalAddress;
  wire       [34:0]   _zz_LsuPlugin_logic_translationStorage_logic_sl_1_write_data_physicalAddress;
  wire       [34:0]   _zz_FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_physicalAddress_1;
  wire       [34:0]   _zz_LsuPlugin_logic_translationStorage_logic_sl_1_write_data_physicalAddress_1;
  wire       [64:0]   _zz_PerformanceCounterPlugin_logic_writePort_data;
  wire       [63:0]   _zz_PerformanceCounterPlugin_logic_counters_cycle_value_2;
  wire       [63:0]   _zz_PerformanceCounterPlugin_logic_counters_instret_value_2;
  wire                decode_ctrls_0_up_isValid;
  wire                fetch_logic_ctrls_0_up_isReady;
  wire                fetch_logic_ctrls_0_up_isValid;
  reg        [63:0]   execute_ctrl5_up_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
  reg                 execute_ctrl5_up_COMMIT_lane0;
  reg        [4:0]    execute_ctrl5_up_RD_PHYS_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_NEED_HIT_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_3_PERM_OK_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_2_PERM_OK_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_1_PERM_OK_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_0_PERM_OK_lane0;
  wire       [11:0]   execute_ctrl3_down_Decode_STORE_ID_lane0;
  wire                execute_ctrl3_down_LsuL1_PREFETCH_lane0;
  wire       [7:0]    execute_ctrl3_down_LsuL1_MASK_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_LSU_PREFETCH_lane0;
  wire                execute_ctrl3_down_AguPlugin_FLOAT_lane0;
  wire                execute_ctrl3_down_AguPlugin_ATOMIC_lane0;
  wire                execute_ctrl3_down_AguPlugin_LOAD_lane0;
  wire                execute_ctrl3_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  wire                execute_ctrl3_down_COMPLETION_AT_4_lane0;
  wire                execute_ctrl3_down_lane0_integer_WriteBackPlugin_SEL_lane0;
  wire                execute_ctrl3_down_MulPlugin_HIGH_lane0;
  wire                execute_ctrl3_down_early0_MulPlugin_SEL_lane0;
  wire       [63:0]   execute_ctrl3_down_integer_RS2_lane0;
  wire       [1:0]    execute_ctrl3_down_AguPlugin_SIZE_lane0;
  wire       [38:0]   execute_ctrl3_down_PC_lane0;
  wire       [0:0]    execute_ctrl3_down_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  wire       [11:0]   execute_ctrl3_down_Prediction_BRANCH_HISTORY_lane0;
  wire       [31:0]   execute_ctrl3_down_Decode_UOP_lane0;
  reg                 execute_ctrl4_up_MMU_BYPASS_TRANSLATION_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_pmpPort_logic_onEntries_3_tor_BIGGER_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_pmpPort_logic_onEntries_3_napot_HIT_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_pmpPort_logic_onEntries_2_tor_BIGGER_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_pmpPort_logic_onEntries_2_napot_HIT_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_pmpPort_logic_onEntries_1_tor_BIGGER_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_pmpPort_logic_onEntries_1_napot_HIT_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_pmpPort_logic_onEntries_0_tor_BIGGER_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_pmpPort_logic_onEntries_0_napot_HIT_lane0;
  reg                 execute_ctrl4_up_MMU_HAZARD_lane0;
  reg                 execute_ctrl4_up_MMU_REFILL_lane0;
  reg                 execute_ctrl4_up_MMU_ACCESS_FAULT_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_MMU_FAILURE_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_MMU_PAGE_FAULT_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_onPma_IO_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_onPma_IO_RSP_lane0_fault;
  reg                 execute_ctrl4_up_LsuPlugin_logic_onPma_IO_RSP_lane0_io;
  reg                 execute_ctrl4_up_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault;
  reg                 execute_ctrl4_up_LsuPlugin_logic_onPma_CACHED_RSP_lane0_io;
  reg                 execute_ctrl4_up_LsuPlugin_logic_preCtrl_IS_AMO_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0;
  reg        [31:0]   execute_ctrl4_up_MMU_TRANSLATED_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_onTrigger_HIT_lane0;
  reg        [25:0]   execute_ctrl4_up_early0_MulPlugin_logic_steps_0_adders_2_lane0;
  reg        [46:0]   execute_ctrl4_up_early0_MulPlugin_logic_steps_0_adders_1_lane0;
  reg        [63:0]   execute_ctrl4_up_early0_MulPlugin_logic_steps_0_adders_0_lane0;
  reg        [1:0]    execute_ctrl4_up_LsuL1Plugin_logic_WAYS_HITS_lane0;
  reg                 execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_loaded;
  reg        [19:0]   execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_address;
  reg                 execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault;
  reg                 execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_loaded;
  reg        [19:0]   execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_address;
  reg                 execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault;
  reg        [31:0]   execute_ctrl4_up_LsuL1_PHYSICAL_ADDRESS_lane0;
  reg        [1:0]    execute_ctrl4_up_LsuL1Plugin_logic_WRITE_TO_READ_HAZARDS_lane0;
  reg        [63:0]   execute_ctrl4_up_LsuL1Plugin_logic_BANKS_MUXES_lane0_0;
  reg        [63:0]   execute_ctrl4_up_LsuL1Plugin_logic_BANKS_MUXES_lane0_1;
  reg        [1:0]    execute_ctrl4_up_LsuL1Plugin_logic_BANK_BUSY_REMAPPED_lane0;
  reg        [0:0]    execute_ctrl4_up_LsuL1Plugin_logic_SHARED_lane0_plru_0;
  reg        [1:0]    execute_ctrl4_up_LsuL1Plugin_logic_SHARED_lane0_dirty;
  reg                 execute_ctrl4_up_LsuPlugin_logic_pmpPort_logic_NEED_HIT_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_pmpPort_logic_onEntries_3_PERM_OK_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_pmpPort_logic_onEntries_2_PERM_OK_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_pmpPort_logic_onEntries_1_PERM_OK_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_pmpPort_logic_onEntries_0_PERM_OK_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_FROM_PREFETCH_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_FROM_LSU_lane0;
  reg        [11:0]   execute_ctrl4_up_Decode_STORE_ID_lane0;
  reg                 execute_ctrl4_up_LsuL1_FLUSH_lane0;
  reg                 execute_ctrl4_up_LsuL1_PREFETCH_lane0;
  reg                 execute_ctrl4_up_LsuL1_INVALID_lane0;
  reg                 execute_ctrl4_up_LsuL1_CLEAN_lane0;
  reg                 execute_ctrl4_up_LsuL1_STORE_lane0;
  reg                 execute_ctrl4_up_LsuL1_ATOMIC_lane0;
  reg                 execute_ctrl4_up_LsuL1_LOAD_lane0;
  reg        [1:0]    execute_ctrl4_up_LsuL1_SIZE_lane0;
  reg        [7:0]    execute_ctrl4_up_LsuL1_MASK_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_FROM_ACCESS_lane0;
  reg        [25:0]   execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_15_lane0;
  reg        [42:0]   execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_14_lane0;
  reg        [42:0]   execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_13_lane0;
  reg        [33:0]   execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_12_lane0;
  reg        [59:0]   execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_11_lane0;
  reg        [59:0]   execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_10_lane0;
  reg        [33:0]   execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_9_lane0;
  reg        [33:0]   execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_8_lane0;
  reg        [76:0]   execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_7_lane0;
  reg        [76:0]   execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_6_lane0;
  reg        [33:0]   execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_5_lane0;
  reg        [33:0]   execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_4_lane0;
  reg        [33:0]   execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_3_lane0;
  reg        [33:0]   execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_2_lane0;
  reg        [33:0]   execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_1_lane0;
  reg        [33:0]   execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_0_lane0;
  reg        [7:0]    execute_ctrl4_up_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0;
  reg        [63:0]   execute_ctrl4_up_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0;
  reg        [38:0]   execute_ctrl4_up_LsuL1_MIXED_ADDRESS_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_LSU_PREFETCH_lane0;
  reg                 execute_ctrl4_up_AguPlugin_FLOAT_lane0;
  reg                 execute_ctrl4_up_AguPlugin_ATOMIC_lane0;
  reg                 execute_ctrl4_up_AguPlugin_STORE_lane0;
  reg                 execute_ctrl4_up_AguPlugin_LOAD_lane0;
  reg        [1:0]    execute_ctrl4_up_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
  reg                 execute_ctrl4_up_lane0_IntFormatPlugin_logic_SIGNED_lane0;
  reg                 execute_ctrl4_up_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  reg                 execute_ctrl4_up_COMPLETION_AT_4_lane0;
  reg                 execute_ctrl4_up_lane0_integer_WriteBackPlugin_SEL_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_FENCE_lane0;
  reg                 execute_ctrl4_up_AguPlugin_SEL_lane0;
  reg                 execute_ctrl4_up_MulPlugin_HIGH_lane0;
  reg                 execute_ctrl4_up_early0_MulPlugin_SEL_lane0;
  reg        [1:0]    execute_ctrl4_up_AguPlugin_SIZE_lane0;
  reg        [4:0]    execute_ctrl4_up_RD_PHYS_lane0;
  reg        [15:0]   execute_ctrl4_up_Decode_UOP_ID_lane0;
  reg        [38:0]   execute_ctrl4_up_PC_lane0;
  reg        [0:0]    execute_ctrl4_up_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  reg        [11:0]   execute_ctrl4_up_Prediction_BRANCH_HISTORY_lane0;
  reg        [31:0]   execute_ctrl4_up_Decode_UOP_lane0;
  wire                execute_ctrl2_down_LsuL1Plugin_logic_FREEZE_HAZARD_lane0;
  wire                execute_ctrl2_down_LsuPlugin_logic_LSU_PREFETCH_lane0;
  wire                execute_ctrl2_down_AguPlugin_FLOAT_lane0;
  wire                execute_ctrl2_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  wire                execute_ctrl2_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  wire                execute_ctrl2_down_COMPLETION_AT_3_lane0;
  wire                execute_ctrl2_down_COMPLETION_AT_4_lane0;
  wire                execute_ctrl2_down_lane0_integer_WriteBackPlugin_SEL_lane0;
  wire                execute_ctrl2_down_MulPlugin_HIGH_lane0;
  wire                execute_ctrl2_down_early0_MulPlugin_SEL_lane0;
  wire       [63:0]   execute_ctrl2_down_integer_RS2_lane0;
  reg        [0:0]    execute_ctrl3_up_MMU_L1_HITS_PRE_VALID_lane0;
  reg                 execute_ctrl3_up_MMU_L1_ENTRIES_lane0_0_valid;
  reg        [12:0]   execute_ctrl3_up_MMU_L1_ENTRIES_lane0_0_virtualAddress;
  reg        [10:0]   execute_ctrl3_up_MMU_L1_ENTRIES_lane0_0_physicalAddress;
  reg                 execute_ctrl3_up_MMU_L1_ENTRIES_lane0_0_allowRead;
  reg                 execute_ctrl3_up_MMU_L1_ENTRIES_lane0_0_allowWrite;
  reg                 execute_ctrl3_up_MMU_L1_ENTRIES_lane0_0_allowExecute;
  reg                 execute_ctrl3_up_MMU_L1_ENTRIES_lane0_0_allowUser;
  reg        [2:0]    execute_ctrl3_up_MMU_L0_HITS_PRE_VALID_lane0;
  reg                 execute_ctrl3_up_MMU_L0_ENTRIES_lane0_0_valid;
  reg        [21:0]   execute_ctrl3_up_MMU_L0_ENTRIES_lane0_0_virtualAddress;
  reg        [19:0]   execute_ctrl3_up_MMU_L0_ENTRIES_lane0_0_physicalAddress;
  reg                 execute_ctrl3_up_MMU_L0_ENTRIES_lane0_0_allowRead;
  reg                 execute_ctrl3_up_MMU_L0_ENTRIES_lane0_0_allowWrite;
  reg                 execute_ctrl3_up_MMU_L0_ENTRIES_lane0_0_allowExecute;
  reg                 execute_ctrl3_up_MMU_L0_ENTRIES_lane0_0_allowUser;
  reg                 execute_ctrl3_up_MMU_L0_ENTRIES_lane0_1_valid;
  reg        [21:0]   execute_ctrl3_up_MMU_L0_ENTRIES_lane0_1_virtualAddress;
  reg        [19:0]   execute_ctrl3_up_MMU_L0_ENTRIES_lane0_1_physicalAddress;
  reg                 execute_ctrl3_up_MMU_L0_ENTRIES_lane0_1_allowRead;
  reg                 execute_ctrl3_up_MMU_L0_ENTRIES_lane0_1_allowWrite;
  reg                 execute_ctrl3_up_MMU_L0_ENTRIES_lane0_1_allowExecute;
  reg                 execute_ctrl3_up_MMU_L0_ENTRIES_lane0_1_allowUser;
  reg                 execute_ctrl3_up_MMU_L0_ENTRIES_lane0_2_valid;
  reg        [21:0]   execute_ctrl3_up_MMU_L0_ENTRIES_lane0_2_virtualAddress;
  reg        [19:0]   execute_ctrl3_up_MMU_L0_ENTRIES_lane0_2_physicalAddress;
  reg                 execute_ctrl3_up_MMU_L0_ENTRIES_lane0_2_allowRead;
  reg                 execute_ctrl3_up_MMU_L0_ENTRIES_lane0_2_allowWrite;
  reg                 execute_ctrl3_up_MMU_L0_ENTRIES_lane0_2_allowExecute;
  reg                 execute_ctrl3_up_MMU_L0_ENTRIES_lane0_2_allowUser;
  reg                 execute_ctrl3_up_LsuPlugin_logic_pmpPort_logic_NEED_HIT_lane0;
  reg                 execute_ctrl3_up_LsuPlugin_logic_pmpPort_logic_onEntries_3_PERM_OK_lane0;
  reg                 execute_ctrl3_up_LsuPlugin_logic_pmpPort_logic_onEntries_2_PERM_OK_lane0;
  reg                 execute_ctrl3_up_LsuPlugin_logic_pmpPort_logic_onEntries_1_PERM_OK_lane0;
  reg                 execute_ctrl3_up_LsuPlugin_logic_pmpPort_logic_onEntries_0_PERM_OK_lane0;
  reg                 execute_ctrl3_up_LsuPlugin_logic_FROM_PREFETCH_lane0;
  reg                 execute_ctrl3_up_LsuPlugin_logic_FROM_LSU_lane0;
  reg        [11:0]   execute_ctrl3_up_Decode_STORE_ID_lane0;
  reg                 execute_ctrl3_up_LsuL1_FLUSH_lane0;
  reg                 execute_ctrl3_up_LsuL1_PREFETCH_lane0;
  reg                 execute_ctrl3_up_LsuL1_INVALID_lane0;
  reg                 execute_ctrl3_up_LsuL1_CLEAN_lane0;
  reg                 execute_ctrl3_up_LsuL1_STORE_lane0;
  reg                 execute_ctrl3_up_LsuL1_ATOMIC_lane0;
  reg                 execute_ctrl3_up_LsuL1_LOAD_lane0;
  reg        [1:0]    execute_ctrl3_up_LsuL1_SIZE_lane0;
  reg        [7:0]    execute_ctrl3_up_LsuL1_MASK_lane0;
  reg                 execute_ctrl3_up_LsuPlugin_logic_FROM_ACCESS_lane0;
  reg                 execute_ctrl3_up_LsuPlugin_logic_FORCE_PHYSICAL_lane0;
  reg        [63:0]   execute_ctrl3_up_DivPlugin_DIV_RESULT_lane0;
  reg        [25:0]   execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_15_lane0;
  reg        [42:0]   execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_14_lane0;
  reg        [42:0]   execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_13_lane0;
  reg        [33:0]   execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_12_lane0;
  reg        [59:0]   execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_11_lane0;
  reg        [59:0]   execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_10_lane0;
  reg        [33:0]   execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_9_lane0;
  reg        [33:0]   execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_8_lane0;
  reg        [76:0]   execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_7_lane0;
  reg        [76:0]   execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_6_lane0;
  reg        [33:0]   execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_5_lane0;
  reg        [33:0]   execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_4_lane0;
  reg        [33:0]   execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_3_lane0;
  reg        [33:0]   execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_2_lane0;
  reg        [33:0]   execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_1_lane0;
  reg        [33:0]   execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_0_lane0;
  reg        [7:0]    execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0;
  reg        [63:0]   execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0;
  reg        [0:0]    execute_ctrl3_up_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_plru_0;
  reg        [1:0]    execute_ctrl3_up_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_dirty;
  reg                 execute_ctrl3_up_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALID_lane0;
  reg        [31:0]   execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_ADDRESS_lane0;
  reg                 execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_VALID_lane0;
  reg        [1:0]    execute_ctrl3_up_LsuL1Plugin_logic_BANK_BUSY_lane0;
  reg        [38:0]   execute_ctrl3_up_LsuL1_MIXED_ADDRESS_lane0;
  reg        [63:0]   execute_ctrl3_up_early0_SrcPlugin_ADD_SUB_lane0;
  reg                 execute_ctrl3_up_COMMIT_lane0;
  reg                 execute_ctrl3_up_LsuPlugin_logic_LSU_PREFETCH_lane0;
  reg                 execute_ctrl3_up_AguPlugin_FLOAT_lane0;
  reg                 execute_ctrl3_up_AguPlugin_ATOMIC_lane0;
  reg                 execute_ctrl3_up_AguPlugin_STORE_lane0;
  reg                 execute_ctrl3_up_AguPlugin_LOAD_lane0;
  reg        [1:0]    execute_ctrl3_up_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
  reg                 execute_ctrl3_up_lane0_IntFormatPlugin_logic_SIGNED_lane0;
  reg                 execute_ctrl3_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  reg                 execute_ctrl3_up_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  reg                 execute_ctrl3_up_COMPLETION_AT_3_lane0;
  reg                 execute_ctrl3_up_COMPLETION_AT_4_lane0;
  reg                 execute_ctrl3_up_lane0_integer_WriteBackPlugin_SEL_lane0;
  reg                 execute_ctrl3_up_LsuPlugin_logic_FENCE_lane0;
  reg                 execute_ctrl3_up_AguPlugin_SEL_lane0;
  reg                 execute_ctrl3_up_CsrAccessPlugin_SEL_lane0;
  reg                 execute_ctrl3_up_MulPlugin_HIGH_lane0;
  reg                 execute_ctrl3_up_early0_DivPlugin_SEL_lane0;
  reg                 execute_ctrl3_up_early0_MulPlugin_SEL_lane0;
  reg        [63:0]   execute_ctrl3_up_integer_RS2_lane0;
  reg        [1:0]    execute_ctrl3_up_AguPlugin_SIZE_lane0;
  reg        [4:0]    execute_ctrl3_up_RD_PHYS_lane0;
  reg        [15:0]   execute_ctrl3_up_Decode_UOP_ID_lane0;
  reg                 execute_ctrl3_up_TRAP_lane0;
  reg        [38:0]   execute_ctrl3_up_PC_lane0;
  reg        [0:0]    execute_ctrl3_up_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  reg        [11:0]   execute_ctrl3_up_Prediction_BRANCH_HISTORY_lane0;
  reg        [31:0]   execute_ctrl3_up_Decode_UOP_lane0;
  wire       [1:0]    execute_ctrl1_down_AguPlugin_SIZE_lane0;
  wire                execute_ctrl1_down_COMPLETED_lane0;
  wire       [4:0]    execute_ctrl1_down_RD_PHYS_lane0;
  wire       [15:0]   execute_ctrl1_down_Decode_UOP_ID_lane0;
  wire       [0:0]    execute_ctrl1_down_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  wire       [11:0]   execute_ctrl1_down_Prediction_BRANCH_HISTORY_lane0;
  wire       [1:0]    execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane0_0;
  wire       [1:0]    execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane0_1;
  wire       [1:0]    execute_ctrl1_down_Prediction_ALIGNED_SLICES_BRANCH_lane0;
  wire       [1:0]    execute_ctrl1_down_Prediction_ALIGNED_SLICES_TAKEN_lane0;
  wire       [38:0]   execute_ctrl1_down_Prediction_ALIGNED_JUMPED_PC_lane0;
  wire                execute_ctrl1_down_Prediction_ALIGNED_JUMPED_lane0;
  wire                execute_ctrl1_down_isReady;
  reg        [2:0]    execute_ctrl2_up_early0_EnvPlugin_OP_lane0;
  reg                 execute_ctrl2_up_LsuPlugin_logic_LSU_PREFETCH_lane0;
  reg                 execute_ctrl2_up_AguPlugin_INVALIDATE_lane0;
  reg                 execute_ctrl2_up_AguPlugin_CLEAN_lane0;
  reg                 execute_ctrl2_up_AguPlugin_FLOAT_lane0;
  reg                 execute_ctrl2_up_AguPlugin_ATOMIC_lane0;
  reg                 execute_ctrl2_up_AguPlugin_STORE_lane0;
  reg                 execute_ctrl2_up_AguPlugin_LOAD_lane0;
  reg                 execute_ctrl2_up_CsrAccessPlugin_CSR_CLEAR_lane0;
  reg                 execute_ctrl2_up_CsrAccessPlugin_CSR_MASK_lane0;
  reg                 execute_ctrl2_up_CsrAccessPlugin_CSR_IMM_lane0;
  reg                 execute_ctrl2_up_RsUnsignedPlugin_IS_W_lane0;
  reg                 execute_ctrl2_up_DivPlugin_REM_lane0;
  reg                 execute_ctrl2_up_RsUnsignedPlugin_RS2_SIGNED_lane0;
  reg                 execute_ctrl2_up_RsUnsignedPlugin_RS1_SIGNED_lane0;
  reg        [1:0]    execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane0;
  reg                 execute_ctrl2_up_BarrelShifterPlugin_IS_W_RIGHT_lane0;
  reg                 execute_ctrl2_up_BarrelShifterPlugin_IS_W_lane0;
  reg                 execute_ctrl2_up_BarrelShifterPlugin_SIGNED_lane0;
  reg                 execute_ctrl2_up_BarrelShifterPlugin_LEFT_lane0;
  reg                 execute_ctrl2_up_SrcStageables_UNSIGNED_lane0;
  reg                 execute_ctrl2_up_BYPASSED_AT_3_lane0;
  reg        [1:0]    execute_ctrl2_up_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
  reg                 execute_ctrl2_up_lane0_IntFormatPlugin_logic_SIGNED_lane0;
  reg                 execute_ctrl2_up_SrcStageables_ZERO_lane0;
  reg                 execute_ctrl2_up_SrcStageables_REVERT_lane0;
  reg        [1:0]    execute_ctrl2_up_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  reg                 execute_ctrl2_up_early0_IntAluPlugin_ALU_SLTX_lane0;
  reg                 execute_ctrl2_up_early0_IntAluPlugin_ALU_ADD_SUB_lane0;
  reg                 execute_ctrl2_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  reg                 execute_ctrl2_up_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  reg                 execute_ctrl2_up_lane0_logic_completions_onCtrl_0_ENABLE_lane0;
  reg                 execute_ctrl2_up_COMPLETION_AT_3_lane0;
  reg                 execute_ctrl2_up_COMPLETION_AT_4_lane0;
  reg                 execute_ctrl2_up_COMPLETION_AT_2_lane0;
  reg                 execute_ctrl2_up_lane0_integer_WriteBackPlugin_SEL_lane0;
  reg                 execute_ctrl2_up_AguPlugin_SEL_lane0;
  reg                 execute_ctrl2_up_CsrAccessPlugin_SEL_lane0;
  reg                 execute_ctrl2_up_MulPlugin_HIGH_lane0;
  reg                 execute_ctrl2_up_early0_EnvPlugin_SEL_lane0;
  reg                 execute_ctrl2_up_early0_DivPlugin_SEL_lane0;
  reg                 execute_ctrl2_up_early0_MulPlugin_SEL_lane0;
  reg                 execute_ctrl2_up_early0_BranchPlugin_SEL_lane0;
  reg                 execute_ctrl2_up_early0_BarrelShifterPlugin_SEL_lane0;
  reg                 execute_ctrl2_up_early0_IntAluPlugin_SEL_lane0;
  reg                 execute_ctrl2_up_MAY_FLUSH_PRECISE_3_lane0;
  reg        [63:0]   execute_ctrl2_up_early0_SrcPlugin_SRC2_lane0;
  reg        [63:0]   execute_ctrl2_up_early0_SrcPlugin_SRC1_lane0;
  reg        [1:0]    execute_ctrl2_up_AguPlugin_SIZE_lane0;
  reg        [15:0]   execute_ctrl2_up_Decode_UOP_ID_lane0;
  reg        [38:0]   execute_ctrl2_up_PC_lane0;
  reg        [0:0]    execute_ctrl2_up_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  reg        [11:0]   execute_ctrl2_up_Prediction_BRANCH_HISTORY_lane0;
  reg        [1:0]    execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane0_0;
  reg        [1:0]    execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane0_1;
  reg        [1:0]    execute_ctrl2_up_Prediction_ALIGNED_SLICES_BRANCH_lane0;
  reg        [1:0]    execute_ctrl2_up_Prediction_ALIGNED_SLICES_TAKEN_lane0;
  reg        [38:0]   execute_ctrl2_up_Prediction_ALIGNED_JUMPED_PC_lane0;
  reg                 execute_ctrl2_up_Prediction_ALIGNED_JUMPED_lane0;
  reg        [31:0]   execute_ctrl2_up_Decode_UOP_lane0;
  wire                execute_ctrl0_down_COMPLETED_lane0;
  wire       [4:0]    execute_ctrl0_down_RD_PHYS_lane0;
  wire                execute_ctrl0_down_TRAP_lane0;
  wire       [38:0]   execute_ctrl0_down_PC_lane0;
  wire       [0:0]    execute_ctrl0_down_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  wire       [11:0]   execute_ctrl0_down_Prediction_BRANCH_HISTORY_lane0;
  wire       [1:0]    execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane0_0;
  wire       [1:0]    execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane0_1;
  wire       [1:0]    execute_ctrl0_down_Prediction_ALIGNED_SLICES_BRANCH_lane0;
  wire       [1:0]    execute_ctrl0_down_Prediction_ALIGNED_SLICES_TAKEN_lane0;
  wire       [38:0]   execute_ctrl0_down_Prediction_ALIGNED_JUMPED_PC_lane0;
  wire                execute_ctrl0_down_Prediction_ALIGNED_JUMPED_lane0;
  reg        [1:0]    execute_ctrl1_up_AguPlugin_SIZE_lane0;
  reg                 execute_ctrl1_up_COMPLETED_lane0;
  reg        [4:0]    execute_ctrl1_up_RS2_PHYS_lane0;
  reg        [4:0]    execute_ctrl1_up_RS1_PHYS_lane0;
  reg        [15:0]   execute_ctrl1_up_Decode_UOP_ID_lane0;
  reg                 execute_ctrl1_up_TRAP_lane0;
  reg        [38:0]   execute_ctrl1_up_PC_lane0;
  reg        [0:0]    execute_ctrl1_up_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  reg        [11:0]   execute_ctrl1_up_Prediction_BRANCH_HISTORY_lane0;
  reg        [1:0]    execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane0_0;
  reg        [1:0]    execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane0_1;
  reg        [1:0]    execute_ctrl1_up_Prediction_ALIGNED_SLICES_BRANCH_lane0;
  reg        [1:0]    execute_ctrl1_up_Prediction_ALIGNED_SLICES_TAKEN_lane0;
  reg        [38:0]   execute_ctrl1_up_Prediction_ALIGNED_JUMPED_PC_lane0;
  reg                 execute_ctrl1_up_Prediction_ALIGNED_JUMPED_lane0;
  reg        [31:0]   execute_ctrl1_up_Decode_UOP_lane0;
  wire                decode_ctrls_1_down_isReady;
  wire                decode_ctrls_0_down_Prediction_ALIGN_REDO_0;
  wire       [1:0]    decode_ctrls_0_down_Prediction_ALIGNED_SLICES_TAKEN_0;
  wire       [1:0]    decode_ctrls_0_down_Prediction_ALIGNED_SLICES_BRANCH_0;
  wire       [38:0]   decode_ctrls_0_down_Prediction_ALIGNED_JUMPED_PC_0;
  wire                decode_ctrls_0_down_Prediction_ALIGNED_JUMPED_0;
  wire       [11:0]   decode_ctrls_0_down_Prediction_BRANCH_HISTORY_0;
  wire       [1:0]    decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_0_0;
  wire       [1:0]    decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_0_1;
  wire       [0:0]    decode_ctrls_0_down_Decode_INSTRUCTION_SLICE_COUNT_0;
  wire       [31:0]   decode_ctrls_0_down_Decode_INSTRUCTION_RAW_0;
  wire                decode_ctrls_0_down_Decode_DECOMPRESSION_FAULT_0;
  wire       [31:0]   decode_ctrls_0_down_Decode_INSTRUCTION_0;
  wire                decode_ctrls_0_down_isValid;
  wire                decode_ctrls_0_down_isReady;
  reg                 decode_ctrls_1_up_Prediction_ALIGN_REDO_0;
  reg        [1:0]    decode_ctrls_1_up_Prediction_ALIGNED_SLICES_TAKEN_0;
  reg        [1:0]    decode_ctrls_1_up_Prediction_ALIGNED_SLICES_BRANCH_0;
  reg        [38:0]   decode_ctrls_1_up_Prediction_ALIGNED_JUMPED_PC_0;
  reg                 decode_ctrls_1_up_Prediction_ALIGNED_JUMPED_0;
  reg        [11:0]   decode_ctrls_1_up_Prediction_BRANCH_HISTORY_0;
  reg        [1:0]    decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_0_0;
  reg        [1:0]    decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_0_1;
  reg        [9:0]    decode_ctrls_1_up_Decode_DOP_ID_0;
  reg        [38:0]   decode_ctrls_1_up_PC_0;
  reg        [0:0]    decode_ctrls_1_up_Decode_INSTRUCTION_SLICE_COUNT_0;
  reg        [31:0]   decode_ctrls_1_up_Decode_INSTRUCTION_RAW_0;
  reg                 decode_ctrls_1_up_Decode_DECOMPRESSION_FAULT_0;
  reg        [31:0]   decode_ctrls_1_up_Decode_INSTRUCTION_0;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_NEED_HIT;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_PERM_OK;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_PERM_OK;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_PERM_OK;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_PERM_OK;
  wire       [9:0]    fetch_logic_ctrls_1_down_Fetch_ID;
  wire                fetch_logic_ctrls_1_down_Fetch_PC_FAULT;
  wire                fetch_logic_ctrls_1_down_isValid;
  wire                fetch_logic_ctrls_1_down_isReady;
  reg                 fetch_logic_ctrls_2_up_MMU_ACCESS_FAULT;
  reg                 fetch_logic_ctrls_2_up_MMU_PAGE_FAULT;
  reg                 fetch_logic_ctrls_2_up_MMU_ALLOW_EXECUTE;
  reg                 fetch_logic_ctrls_2_up_MMU_REFILL;
  reg                 fetch_logic_ctrls_2_up_MMU_HAZARD;
  reg        [1:0]    fetch_logic_ctrls_2_up_Prediction_WORD_SLICES_TAKEN;
  reg        [1:0]    fetch_logic_ctrls_2_up_Prediction_WORD_SLICES_BRANCH;
  reg        [38:0]   fetch_logic_ctrls_2_up_Prediction_WORD_JUMP_PC;
  reg        [0:0]    fetch_logic_ctrls_2_up_Prediction_WORD_JUMP_SLICE;
  reg                 fetch_logic_ctrls_2_up_Prediction_WORD_JUMPED;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_tor_BIGGER;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_napot_HIT;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_tor_BIGGER;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_napot_HIT;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_tor_BIGGER;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_napot_HIT;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_tor_BIGGER;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_napot_HIT;
  reg        [31:0]   fetch_logic_ctrls_2_up_MMU_TRANSLATED;
  reg        [1:0]    fetch_logic_ctrls_2_up_GSharePlugin_GSHARE_COUNTER_0;
  reg        [1:0]    fetch_logic_ctrls_2_up_GSharePlugin_GSHARE_COUNTER_1;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_HIT;
  reg                 fetch_logic_ctrls_2_up_MMU_BYPASS_TRANSLATION;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_HITS_0;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_HITS_1;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_HAZARD;
  reg        [31:0]   fetch_logic_ctrls_2_up_FetchL1Plugin_logic_BANKS_MUXES_0;
  reg        [31:0]   fetch_logic_ctrls_2_up_FetchL1Plugin_logic_BANKS_MUXES_1;
  reg        [0:0]    fetch_logic_ctrls_2_up_FetchL1Plugin_logic_PLRU_BYPASSED_0;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_0_loaded;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_0_error;
  reg        [19:0]   fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_0_address;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_1_loaded;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_1_error;
  reg        [19:0]   fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_1_address;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_pmpPort_logic_NEED_HIT;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_PERM_OK;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_PERM_OK;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_PERM_OK;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_PERM_OK;
  reg        [11:0]   fetch_logic_ctrls_2_up_Prediction_BRANCH_HISTORY;
  reg        [9:0]    fetch_logic_ctrls_2_up_Fetch_ID;
  reg                 fetch_logic_ctrls_2_up_Fetch_PC_FAULT;
  reg        [38:0]   fetch_logic_ctrls_2_up_Fetch_WORD_PC;
  wire                fetch_logic_ctrls_0_down_Fetch_PC_FAULT;
  wire                fetch_logic_ctrls_0_down_isValid;
  reg        [0:0]    fetch_logic_ctrls_1_up_BtbPlugin_logic_readCmd_HAZARDS;
  reg                 fetch_logic_ctrls_1_up_FetchL1Plugin_logic_pmpPort_logic_NEED_HIT;
  reg                 fetch_logic_ctrls_1_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_PERM_OK;
  reg                 fetch_logic_ctrls_1_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_PERM_OK;
  reg                 fetch_logic_ctrls_1_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_PERM_OK;
  reg                 fetch_logic_ctrls_1_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_PERM_OK;
  reg                 fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_valid;
  reg        [12:0]   fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_address;
  reg        [1:0]    fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_data_0;
  reg        [1:0]    fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_data_1;
  reg        [11:0]   fetch_logic_ctrls_1_up_Prediction_BRANCH_HISTORY;
  reg        [12:0]   fetch_logic_ctrls_1_up_GSharePlugin_logic_HASH;
  reg        [5:0]    fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_TAGS_UPDATE_ADDRESS;
  reg                 fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_TAGS_UPDATE;
  reg        [0:0]    fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_0;
  reg                 fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_PLRU_BYPASS_VALID;
  reg                 _zz_1;
  reg        [9:0]    fetch_logic_ctrls_1_up_Fetch_ID;
  reg                 fetch_logic_ctrls_1_up_Fetch_PC_FAULT;
  reg        [38:0]   fetch_logic_ctrls_1_up_Fetch_WORD_PC;
  reg                 fetch_logic_ctrls_2_up_valid;
  wire                decode_ctrls_1_down_valid;
  reg                 fetch_logic_ctrls_1_down_valid;
  wire                decode_ctrls_0_down_valid;
  reg                 fetch_logic_ctrls_0_down_valid;
  wire                execute_ctrl0_up_ready;
  wire                execute_ctrl0_down_ready;
  wire                execute_ctrl1_up_ready;
  wire                execute_ctrl1_down_ready;
  wire                execute_ctrl2_up_ready;
  wire                execute_ctrl2_down_ready;
  wire                execute_ctrl3_up_ready;
  wire                execute_ctrl3_down_ready;
  wire                fetch_logic_ctrls_0_down_ready;
  wire                execute_ctrl4_up_ready;
  wire                decode_ctrls_0_up_ready;
  wire                fetch_logic_ctrls_1_up_cancel;
  wire                execute_ctrl4_down_ready;
  reg                 decode_ctrls_0_down_ready;
  wire                fetch_logic_ctrls_1_down_ready;
  wire                execute_ctrl5_up_ready;
  wire                fetch_logic_ctrls_2_up_ready;
  wire                fetch_logic_ctrls_2_up_cancel;
  wire                execute_ctrl5_down_ready;
  wire                execute_ctrl4_down_AguPlugin_ATOMIC_lane0;
  wire       [11:0]   execute_ctrl4_down_Decode_STORE_ID_lane0;
  wire       [31:0]   execute_ctrl4_down_MMU_TRANSLATED_lane0;
  wire       [1:0]    execute_ctrl4_down_AguPlugin_SIZE_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_LSU_PREFETCH_lane0;
  wire                execute_ctrl4_down_AguPlugin_LOAD_lane0;
  wire                execute_ctrl4_down_RD_ENABLE_lane0;
  reg                 execute_ctrl4_RD_ENABLE_lane0_bypass;
  reg                 execute_ctrl4_LANE_SEL_lane0_bypass;
  wire                execute_ctrl3_down_RD_ENABLE_lane0;
  reg                 execute_ctrl3_RD_ENABLE_lane0_bypass;
  reg                 execute_ctrl3_LANE_SEL_lane0_bypass;
  wire                execute_ctrl2_down_RD_ENABLE_lane0;
  reg                 execute_ctrl2_RD_ENABLE_lane0_bypass;
  reg                 execute_ctrl2_LANE_SEL_lane0_bypass;
  wire                execute_ctrl1_down_RD_ENABLE_lane0;
  reg                 execute_ctrl1_RD_ENABLE_lane0_bypass;
  wire                execute_ctrl1_down_LANE_SEL_lane0;
  reg                 execute_ctrl1_LANE_SEL_lane0_bypass;
  wire                execute_ctrl0_down_RD_ENABLE_lane0;
  reg                 execute_ctrl0_RD_ENABLE_lane0_bypass;
  reg                 execute_ctrl0_LANE_SEL_lane0_bypass;
  wire                execute_ctrl1_down_TRAP_lane0;
  wire       [2:0]    execute_ctrl1_down_early0_EnvPlugin_OP_lane0;
  wire                execute_ctrl1_down_LsuPlugin_logic_LSU_PREFETCH_lane0;
  wire                execute_ctrl1_down_AguPlugin_INVALIDATE_lane0;
  wire                execute_ctrl1_down_AguPlugin_CLEAN_lane0;
  wire                execute_ctrl1_down_AguPlugin_FLOAT_lane0;
  wire                execute_ctrl1_down_AguPlugin_ATOMIC_lane0;
  wire                execute_ctrl1_down_AguPlugin_STORE_lane0;
  wire                execute_ctrl1_down_AguPlugin_LOAD_lane0;
  wire                execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0;
  wire                execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0;
  wire                execute_ctrl1_down_CsrAccessPlugin_CSR_IMM_lane0;
  wire                execute_ctrl1_down_RsUnsignedPlugin_IS_W_lane0;
  wire                execute_ctrl1_down_DivPlugin_REM_lane0;
  wire                execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0;
  wire                execute_ctrl1_down_RsUnsignedPlugin_RS1_SIGNED_lane0;
  wire       [1:0]    execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0;
  wire                execute_ctrl1_down_BarrelShifterPlugin_IS_W_RIGHT_lane0;
  wire                execute_ctrl1_down_BarrelShifterPlugin_IS_W_lane0;
  wire                execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane0;
  wire                execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0;
  wire                execute_ctrl1_down_SrcStageables_UNSIGNED_lane0;
  wire                execute_ctrl1_down_BYPASSED_AT_3_lane0;
  wire       [1:0]    execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
  wire                execute_ctrl1_down_lane0_IntFormatPlugin_logic_SIGNED_lane0;
  wire                execute_ctrl1_down_SrcStageables_ZERO_lane0;
  wire                execute_ctrl1_down_SrcStageables_REVERT_lane0;
  wire       [1:0]    execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  wire                execute_ctrl1_down_early0_IntAluPlugin_ALU_SLTX_lane0;
  wire                execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0;
  reg                 execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  reg                 execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  reg                 execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0;
  reg                 execute_ctrl1_down_COMPLETION_AT_3_lane0;
  reg                 execute_ctrl1_down_COMPLETION_AT_4_lane0;
  reg                 execute_ctrl1_down_COMPLETION_AT_2_lane0;
  reg                 execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0;
  reg                 execute_ctrl1_down_LsuPlugin_logic_FENCE_lane0;
  reg                 execute_ctrl1_down_AguPlugin_SEL_lane0;
  reg                 execute_ctrl1_down_CsrAccessPlugin_SEL_lane0;
  reg                 execute_ctrl1_down_MulPlugin_HIGH_lane0;
  reg                 execute_ctrl1_down_early0_EnvPlugin_SEL_lane0;
  reg                 execute_ctrl1_down_early0_DivPlugin_SEL_lane0;
  reg                 execute_ctrl1_down_early0_MulPlugin_SEL_lane0;
  reg                 execute_ctrl1_down_early0_BranchPlugin_SEL_lane0;
  reg                 execute_ctrl1_down_early0_BarrelShifterPlugin_SEL_lane0;
  reg                 execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0;
  wire                execute_ctrl3_down_TRAP_lane0;
  wire                execute_ctrl3_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  wire                execute_ctrl4_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  wire                execute_ctrl2_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0;
  wire       [4:0]    execute_ctrl1_down_RS2_PHYS_lane0;
  wire       [4:0]    execute_ctrl0_down_RS2_PHYS_lane0;
  wire       [63:0]   execute_ctrl5_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
  wire       [4:0]    execute_ctrl5_down_RD_PHYS_lane0;
  reg                 execute_ctrl5_up_RD_ENABLE_lane0;
  reg                 execute_ctrl5_up_LANE_SEL_lane0;
  wire       [4:0]    execute_ctrl3_down_RD_PHYS_lane0;
  wire       [4:0]    execute_ctrl1_down_RS1_PHYS_lane0;
  wire       [4:0]    execute_ctrl0_down_RS1_PHYS_lane0;
  reg                 _zz_2;
  wire                execute_ctrl3_down_CsrAccessPlugin_SEL_lane0;
  wire       [4:0]    execute_ctrl2_down_RD_PHYS_lane0;
  wire                execute_ctrl2_down_CsrAccessPlugin_CSR_CLEAR_lane0;
  wire                execute_ctrl2_down_CsrAccessPlugin_CSR_MASK_lane0;
  wire                execute_ctrl2_down_CsrAccessPlugin_CSR_IMM_lane0;
  wire                execute_ctrl2_down_CsrAccessPlugin_SEL_lane0;
  reg                 fetch_logic_ctrls_1_down_MMU_ACCESS_FAULT;
  reg                 fetch_logic_ctrls_1_down_MMU_PAGE_FAULT;
  reg                 fetch_logic_ctrls_1_down_MMU_ALLOW_WRITE;
  reg                 fetch_logic_ctrls_1_down_MMU_ALLOW_READ;
  reg                 fetch_logic_ctrls_1_down_MMU_ALLOW_EXECUTE;
  reg                 fetch_logic_ctrls_1_down_MMU_REFILL;
  reg                 fetch_logic_ctrls_1_down_MMU_HAZARD;
  wire       [0:0]    fetch_logic_ctrls_1_down_MMU_L1_HITS;
  wire       [0:0]    fetch_logic_ctrls_1_down_MMU_L1_HITS_PRE_VALID;
  wire                fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_valid;
  wire       [12:0]   fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_virtualAddress;
  wire       [10:0]   fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_physicalAddress;
  wire                fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_allowRead;
  wire                fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_allowWrite;
  wire                fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_allowExecute;
  wire                fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_allowUser;
  reg        [1:0]    fetch_logic_ctrls_1_down_MMU_L0_HITS;
  reg        [1:0]    fetch_logic_ctrls_1_down_MMU_L0_HITS_PRE_VALID;
  wire                fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_valid;
  wire       [21:0]   fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_virtualAddress;
  wire       [19:0]   fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_physicalAddress;
  wire                fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_allowRead;
  wire                fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_allowWrite;
  wire                fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_allowExecute;
  wire                fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_allowUser;
  wire                fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_valid;
  wire       [21:0]   fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_virtualAddress;
  wire       [19:0]   fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_physicalAddress;
  wire                fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_allowRead;
  wire                fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_allowWrite;
  wire                fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_allowExecute;
  wire                fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_allowUser;
  wire       [31:0]   execute_ctrl3_down_MMU_WAYS_PHYSICAL_lane0_0;
  wire       [31:0]   execute_ctrl3_down_MMU_WAYS_PHYSICAL_lane0_1;
  wire       [31:0]   execute_ctrl3_down_MMU_WAYS_PHYSICAL_lane0_2;
  wire       [31:0]   execute_ctrl3_down_MMU_WAYS_PHYSICAL_lane0_3;
  wire       [3:0]    execute_ctrl3_down_MMU_WAYS_OH_lane0;
  wire                execute_ctrl3_down_MMU_BYPASS_TRANSLATION_lane0;
  reg                 execute_ctrl3_down_MMU_ALLOW_EXECUTE_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_FORCE_PHYSICAL_lane0;
  wire                execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_valid;
  wire       [12:0]   execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_virtualAddress;
  wire       [10:0]   execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_physicalAddress;
  wire                execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_allowRead;
  wire                execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_allowWrite;
  wire                execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_allowExecute;
  wire                execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_allowUser;
  wire       [0:0]    execute_ctrl3_down_MMU_L1_HITS_PRE_VALID_lane0;
  wire       [0:0]    execute_ctrl3_down_MMU_L1_HITS_lane0;
  wire       [0:0]    execute_ctrl2_down_MMU_L1_HITS_PRE_VALID_lane0;
  wire                execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_valid;
  wire       [12:0]   execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_virtualAddress;
  wire       [10:0]   execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_physicalAddress;
  wire                execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_allowRead;
  wire                execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_allowWrite;
  wire                execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_allowExecute;
  wire                execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_allowUser;
  wire                execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_valid;
  wire       [21:0]   execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_virtualAddress;
  wire       [19:0]   execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_physicalAddress;
  wire                execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_allowRead;
  wire                execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_allowWrite;
  wire                execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_allowExecute;
  wire                execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_allowUser;
  wire                execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_valid;
  wire       [21:0]   execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_virtualAddress;
  wire       [19:0]   execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_physicalAddress;
  wire                execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_allowRead;
  wire                execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_allowWrite;
  wire                execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_allowExecute;
  wire                execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_allowUser;
  wire                execute_ctrl3_down_MMU_L0_ENTRIES_lane0_2_valid;
  wire       [21:0]   execute_ctrl3_down_MMU_L0_ENTRIES_lane0_2_virtualAddress;
  wire       [19:0]   execute_ctrl3_down_MMU_L0_ENTRIES_lane0_2_physicalAddress;
  wire                execute_ctrl3_down_MMU_L0_ENTRIES_lane0_2_allowRead;
  wire                execute_ctrl3_down_MMU_L0_ENTRIES_lane0_2_allowWrite;
  wire                execute_ctrl3_down_MMU_L0_ENTRIES_lane0_2_allowExecute;
  wire                execute_ctrl3_down_MMU_L0_ENTRIES_lane0_2_allowUser;
  wire       [2:0]    execute_ctrl3_down_MMU_L0_HITS_PRE_VALID_lane0;
  reg        [2:0]    execute_ctrl3_down_MMU_L0_HITS_lane0;
  reg        [2:0]    execute_ctrl2_down_MMU_L0_HITS_PRE_VALID_lane0;
  wire                execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_valid;
  wire       [21:0]   execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_virtualAddress;
  wire       [19:0]   execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_physicalAddress;
  wire                execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_allowRead;
  wire                execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_allowWrite;
  wire                execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_allowExecute;
  wire                execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_allowUser;
  wire                execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_valid;
  wire       [21:0]   execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_virtualAddress;
  wire       [19:0]   execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_physicalAddress;
  wire                execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_allowRead;
  wire                execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_allowWrite;
  wire                execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_allowExecute;
  wire                execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_allowUser;
  wire                execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_valid;
  wire       [21:0]   execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_virtualAddress;
  wire       [19:0]   execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_physicalAddress;
  wire                execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_allowRead;
  wire                execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_allowWrite;
  wire                execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_allowExecute;
  wire                execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_allowUser;
  wire                fetch_logic_ctrls_0_up_isFiring;
  reg        [9:0]    fetch_logic_ctrls_0_up_Fetch_ID;
  wire                fetch_logic_ctrls_0_up_Fetch_PC_FAULT;
  wire       [38:0]   fetch_logic_ctrls_0_up_Fetch_WORD_PC;
  reg                 fetch_logic_ctrls_0_up_ready;
  wire                fetch_logic_ctrls_0_up_valid;
  reg                 PcPlugin_logic_harts_0_aggregator_fault_1;
  reg        [38:0]   PcPlugin_logic_harts_0_aggregator_target_1;
  wire       [0:0]    execute_ctrl4_down_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  wire       [11:0]   execute_ctrl4_down_Prediction_BRANCH_HISTORY_lane0;
  wire                execute_ctrl5_down_COMMIT_lane0;
  wire                execute_ctrl5_down_isReady;
  wire                execute_ctrl5_down_LANE_SEL_lane0;
  wire                decode_ctrls_0_down_TRAP_0;
  wire                decode_ctrls_1_down_LANE_SEL_0;
  reg                 decode_ctrls_1_LANE_SEL_0_bypass;
  wire                decode_ctrls_0_down_LANE_SEL_0;
  reg                 decode_ctrls_0_LANE_SEL_0_bypass;
  wire                decode_ctrls_0_up_isMoving;
  reg        [1:0]    fetch_logic_ctrls_1_down_Prediction_WORD_SLICES_TAKEN;
  reg        [1:0]    fetch_logic_ctrls_1_down_Prediction_WORD_SLICES_BRANCH;
  wire       [11:0]   fetch_logic_ctrls_1_down_Prediction_BRANCH_HISTORY;
  wire       [38:0]   fetch_logic_ctrls_1_down_Prediction_WORD_JUMP_PC;
  wire       [0:0]    fetch_logic_ctrls_1_down_Prediction_WORD_JUMP_SLICE;
  wire                fetch_logic_ctrls_1_down_Prediction_WORD_JUMPED;
  wire                fetch_logic_ctrls_1_up_isCancel;
  wire                fetch_logic_ctrls_1_up_isReady;
  wire                fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_predict_TAKEN;
  wire       [0:0]    fetch_logic_ctrls_1_down_BtbPlugin_logic_readCmd_HAZARDS;
  wire                fetch_logic_ctrls_1_up_isValid;
  wire                fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_hitCalc_HIT;
  (* keep , syn_keep *) wire       [15:0]   fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_hash /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [0:0]    fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_sliceLow /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [37:0]   fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_pcTarget /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isBranch /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isPush /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isPop /* synthesis syn_keep = 1 */ ;
  wire       [0:0]    fetch_logic_ctrls_0_down_BtbPlugin_logic_readCmd_HAZARDS;
  wire       [15:0]   execute_ctrl0_down_Decode_UOP_ID_lane0;
  wire                execute_ctrl0_down_isReady;
  wire                execute_ctrl0_down_LANE_SEL_lane0;
  wire       [9:0]    decode_ctrls_1_down_Decode_DOP_ID_0;
  wire                decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_0;
  wire                decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_0;
  wire       [4:0]    execute_ctrl4_down_RD_PHYS_lane0;
  wire                execute_ctrl4_down_lane0_integer_WriteBackPlugin_SEL_lane0;
  reg                 execute_ctrl4_up_RD_ENABLE_lane0;
  wire       [63:0]   execute_ctrl4_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
  wire       [63:0]   execute_ctrl4_lane0_integer_WriteBackPlugin_logic_DATA_lane0_bypass;
  reg        [63:0]   execute_ctrl4_up_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
  wire       [15:0]   execute_ctrl3_down_Decode_UOP_ID_lane0;
  wire                execute_ctrl3_down_COMMIT_lane0;
  reg                 execute_ctrl3_up_RD_ENABLE_lane0;
  wire                execute_ctrl3_down_isReady;
  wire                execute_ctrl3_down_LANE_SEL_lane0;
  wire       [63:0]   execute_ctrl3_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
  wire       [63:0]   execute_ctrl3_lane0_integer_WriteBackPlugin_logic_DATA_lane0_bypass;
  reg        [63:0]   execute_ctrl3_up_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
  wire                execute_ctrl2_down_LANE_SEL_lane0;
  wire       [63:0]   execute_ctrl2_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
  wire       [63:0]   execute_ctrl2_lane0_integer_WriteBackPlugin_logic_DATA_lane0_bypass;
  wire                execute_ctrl0_up_COMPLETED_lane0;
  wire                execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_lane0;
  wire                execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_lane0;
  wire       [4:0]    execute_ctrl0_up_RD_PHYS_lane0;
  reg                 execute_ctrl0_up_RD_ENABLE_lane0;
  wire       [4:0]    execute_ctrl0_up_RS2_PHYS_lane0;
  wire                execute_ctrl0_up_RS2_ENABLE_lane0;
  wire       [4:0]    execute_ctrl0_up_RS1_PHYS_lane0;
  wire                execute_ctrl0_up_RS1_ENABLE_lane0;
  wire       [15:0]   execute_ctrl0_up_Decode_UOP_ID_lane0;
  wire                execute_ctrl0_up_TRAP_lane0;
  wire       [38:0]   execute_ctrl0_up_PC_lane0;
  wire                execute_ctrl0_up_DONT_FLUSH_PRECISE_4_lane0;
  wire                execute_ctrl0_up_DONT_FLUSH_PRECISE_3_lane0;
  wire       [0:0]    execute_ctrl0_up_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  wire                execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_FROM_LANES_lane0;
  wire                execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_lane0;
  reg                 execute_ctrl0_up_DispatchPlugin_MAY_FLUSH_lane0;
  wire                execute_ctrl0_up_DispatchPlugin_FENCE_OLDER_lane0;
  wire       [11:0]   execute_ctrl0_up_Prediction_BRANCH_HISTORY_lane0;
  wire       [1:0]    execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0;
  wire       [1:0]    execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_1;
  wire       [1:0]    execute_ctrl0_up_Prediction_ALIGNED_SLICES_BRANCH_lane0;
  wire       [1:0]    execute_ctrl0_up_Prediction_ALIGNED_SLICES_TAKEN_lane0;
  wire       [38:0]   execute_ctrl0_up_Prediction_ALIGNED_JUMPED_PC_lane0;
  wire                execute_ctrl0_up_Prediction_ALIGNED_JUMPED_lane0;
  wire       [31:0]   execute_ctrl0_up_Decode_UOP_lane0;
  wire                execute_ctrl0_up_LANE_SEL_lane0;
  wire                decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0;
  wire                decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_0;
  wire                decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0;
  wire                decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_0;
  wire                decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_0;
  wire                decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_0;
  wire                decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_0;
  wire                decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_0;
  wire       [11:0]   decode_ctrls_1_down_Prediction_BRANCH_HISTORY_0;
  wire       [1:0]    decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0_0;
  wire       [1:0]    decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0_1;
  wire       [1:0]    decode_ctrls_1_down_Prediction_ALIGNED_SLICES_BRANCH_0;
  wire       [1:0]    decode_ctrls_1_down_Prediction_ALIGNED_SLICES_TAKEN_0;
  wire       [38:0]   decode_ctrls_1_down_Prediction_ALIGNED_JUMPED_PC_0;
  wire                decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0;
  wire                decode_ctrls_1_up_isValid;
  reg                 decode_ctrls_1_down_ready;
  wire                execute_ctrl2_down_MAY_FLUSH_PRECISE_3_lane0;
  wire                execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane0;
  wire                execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane0;
  wire                execute_ctrl2_down_BYPASSED_AT_3_lane0;
  reg        [4:0]    execute_ctrl2_up_RD_PHYS_lane0;
  reg                 execute_ctrl2_up_RD_ENABLE_lane0;
  wire                execute_ctrl1_down_BYPASSED_AT_2_lane0;
  reg        [4:0]    execute_ctrl1_up_RD_PHYS_lane0;
  reg                 execute_ctrl1_up_RD_ENABLE_lane0;
  wire       [31:0]   decode_ctrls_1_down_Decode_UOP_0;
  reg                 decode_ctrls_1_up_TRAP_0;
  reg                 decode_ctrls_1_TRAP_0_bypass;
  wire       [15:0]   decode_ctrls_1_down_Decode_UOP_ID_0;
  wire                decode_ctrls_1_up_isReady;
  wire                decode_ctrls_1_down_TRAP_0;
  wire       [0:0]    decode_ctrls_1_down_Decode_INSTRUCTION_SLICE_COUNT_0;
  wire       [38:0]   decode_ctrls_1_down_PC_0;
  wire                decode_ctrls_1_down_Prediction_ALIGN_REDO_0;
  wire                decode_ctrls_1_down_Prediction_ALIGNED_JUMPED_0;
  reg                 decode_ctrls_1_up_LANE_SEL_0;
  wire       [31:0]   decode_ctrls_1_down_Decode_INSTRUCTION_RAW_0;
  wire                decode_ctrls_1_down_AguPlugin_CLEAN_0;
  wire                decode_ctrls_1_down_AguPlugin_INVALIDATE_0;
  wire                decode_ctrls_1_down_Decode_DECOMPRESSION_FAULT_0;
  reg                 decode_ctrls_1_down_Decode_LEGAL_0;
  wire       [4:0]    decode_ctrls_1_down_RD_PHYS_0;
  reg                 decode_ctrls_1_down_RD_ENABLE_0;
  wire       [4:0]    decode_ctrls_1_down_RS2_PHYS_0;
  wire                decode_ctrls_1_down_RS2_ENABLE_0;
  wire       [4:0]    decode_ctrls_1_down_RS1_PHYS_0;
  wire       [31:0]   decode_ctrls_1_down_Decode_INSTRUCTION_0;
  wire                decode_ctrls_1_down_RS1_ENABLE_0;
  wire                decode_ctrls_1_up_isCanceling;
  wire                decode_ctrls_1_up_ready;
  reg                 decode_ctrls_1_up_valid;
  wire                decode_ctrls_1_up_isMoving;
  wire                execute_ctrl3_down_COMPLETION_AT_3_lane0;
  reg                 execute_ctrl3_up_COMPLETED_lane0;
  wire                execute_ctrl3_down_COMPLETED_lane0;
  wire                execute_ctrl3_COMPLETED_lane0_bypass;
  wire                execute_ctrl4_down_COMPLETION_AT_4_lane0;
  reg                 execute_ctrl4_up_COMPLETED_lane0;
  wire                execute_ctrl4_down_COMPLETED_lane0;
  wire                execute_ctrl4_COMPLETED_lane0_bypass;
  wire                execute_ctrl2_down_COMPLETION_AT_2_lane0;
  reg                 execute_ctrl2_up_COMPLETED_lane0;
  wire                execute_ctrl2_down_COMPLETED_lane0;
  wire                execute_ctrl2_COMPLETED_lane0_bypass;
  reg                 execute_ctrl1_up_LANE_SEL_lane0;
  wire       [1:0]    execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane0_0;
  wire       [1:0]    execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane0_1;
  wire                execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_IS_JALR_lane0;
  wire                execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_IS_JAL_lane0;
  wire                execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_MISSALIGNED_lane0;
  reg        [11:0]   early0_BranchPlugin_logic_jumpLogic_history_shifter_2;
  reg        [11:0]   early0_BranchPlugin_logic_jumpLogic_history_shifter_1;
  wire       [1:0]    execute_ctrl2_down_Prediction_ALIGNED_SLICES_TAKEN_lane0;
  wire       [1:0]    execute_ctrl2_down_Prediction_ALIGNED_SLICES_BRANCH_lane0;
  wire       [11:0]   execute_ctrl2_down_Prediction_BRANCH_HISTORY_lane0;
  wire                execute_ctrl2_down_early0_BranchPlugin_SEL_lane0;
  wire                execute_ctrl2_down_Prediction_ALIGNED_JUMPED_lane0;
  wire       [38:0]   execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_btb_REAL_TARGET_lane0;
  wire                execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0;
  wire                execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0;
  wire                execute_ctrl2_down_early0_BranchPlugin_logic_alu_btb_BAD_TARGET_lane0;
  wire       [38:0]   execute_ctrl2_down_Prediction_ALIGNED_JUMPED_PC_lane0;
  wire                execute_ctrl2_down_early0_BranchPlugin_logic_alu_EQ_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_3_PERM_OK_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_2_PERM_OK_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_1_PERM_OK_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_0_PERM_OK_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_NEED_HIT_lane0;
  wire                execute_ctrl2_down_LsuPlugin_logic_pmpPort_logic_NEED_HIT_lane0;
  wire                execute_ctrl2_down_LsuPlugin_logic_pmpPort_logic_onEntries_3_PERM_OK_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_3_HIT_ANY_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_3_napot_HIT_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_3_tor_HIT_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_3_tor_BIGGER_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_3_tor_BIGGER_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_3_napot_HIT_lane0;
  wire       [19:0]   execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_3_napot_MATCH_lane0;
  wire                execute_ctrl2_down_LsuPlugin_logic_pmpPort_logic_onEntries_2_PERM_OK_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_2_HIT_ANY_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_2_napot_HIT_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_2_tor_HIT_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_2_tor_BIGGER_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_2_tor_BIGGER_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_2_napot_HIT_lane0;
  wire       [19:0]   execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_2_napot_MATCH_lane0;
  wire                execute_ctrl2_down_LsuPlugin_logic_pmpPort_logic_onEntries_1_PERM_OK_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_1_HIT_ANY_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_1_napot_HIT_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_1_tor_HIT_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_1_tor_BIGGER_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_1_tor_BIGGER_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_1_napot_HIT_lane0;
  wire       [19:0]   execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_1_napot_MATCH_lane0;
  wire                execute_ctrl2_down_LsuPlugin_logic_pmpPort_logic_onEntries_0_PERM_OK_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_0_HIT_ANY_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_0_napot_HIT_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_0_tor_HIT_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_0_tor_BIGGER_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_0_tor_BIGGER_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_0_napot_HIT_lane0;
  wire       [19:0]   execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_0_napot_MATCH_lane0;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_PERM_OK;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_PERM_OK;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_PERM_OK;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_PERM_OK;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_NEED_HIT;
  wire                fetch_logic_ctrls_0_down_FetchL1Plugin_logic_pmpPort_logic_NEED_HIT;
  wire                fetch_logic_ctrls_0_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_PERM_OK;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_HIT_ANY;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_napot_HIT;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_tor_HIT;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_tor_BIGGER;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_tor_BIGGER;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_napot_HIT;
  wire       [19:0]   fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_napot_MATCH;
  wire                fetch_logic_ctrls_0_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_PERM_OK;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_HIT_ANY;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_napot_HIT;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_tor_HIT;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_tor_BIGGER;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_tor_BIGGER;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_napot_HIT;
  wire       [19:0]   fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_napot_MATCH;
  wire                fetch_logic_ctrls_0_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_PERM_OK;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_HIT_ANY;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_napot_HIT;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_tor_HIT;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_tor_BIGGER;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_tor_BIGGER;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_napot_HIT;
  wire       [19:0]   fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_napot_MATCH;
  wire                fetch_logic_ctrls_0_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_PERM_OK;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_HIT_ANY;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_napot_HIT;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_tor_HIT;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_tor_BIGGER;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_tor_BIGGER;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_napot_HIT;
  wire       [19:0]   fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_napot_MATCH;
  reg        [31:0]   fetch_logic_ctrls_1_down_MMU_TRANSLATED;
  wire                execute_ctrl2_up_COMMIT_lane0;
  wire                execute_ctrl2_down_COMMIT_lane0;
  reg                 execute_ctrl2_COMMIT_lane0_bypass;
  reg                 execute_ctrl2_up_TRAP_lane0;
  wire                execute_ctrl2_down_TRAP_lane0;
  reg                 execute_ctrl2_TRAP_lane0_bypass;
  wire                execute_ctrl2_down_early0_EnvPlugin_SEL_lane0;
  wire       [38:0]   fetch_logic_ctrls_2_down_Prediction_WORD_JUMP_PC;
  wire       [1:0]    fetch_logic_ctrls_2_down_Prediction_WORD_SLICES_TAKEN;
  wire       [1:0]    fetch_logic_ctrls_2_down_Prediction_WORD_SLICES_BRANCH;
  wire       [11:0]   fetch_logic_ctrls_2_down_Prediction_BRANCH_HISTORY;
  wire       [1:0]    fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_1;
  wire       [9:0]    fetch_logic_ctrls_2_down_Fetch_ID;
  wire                fetch_logic_ctrls_2_down_isCancel;
  wire                fetch_logic_ctrls_2_down_ready;
  wire                decode_ctrls_0_up_isCancel;
  wire                fetch_logic_ctrls_2_down_valid;
  wire                fetch_logic_ctrls_2_down_isValid;
  wire                decode_ctrls_0_up_valid;
  wire                decode_ctrls_0_up_Prediction_ALIGN_REDO_0;
  wire       [1:0]    decode_ctrls_0_up_Prediction_ALIGNED_SLICES_TAKEN_0;
  wire       [1:0]    decode_ctrls_0_up_Prediction_ALIGNED_SLICES_BRANCH_0;
  wire       [38:0]   decode_ctrls_0_up_Prediction_ALIGNED_JUMPED_PC_0;
  wire                decode_ctrls_0_up_Prediction_ALIGNED_JUMPED_0;
  wire                decode_ctrls_0_up_TRAP_0;
  wire       [0:0]    decode_ctrls_0_up_Prediction_WORD_JUMP_SLICE_0;
  wire                decode_ctrls_0_up_Prediction_WORD_JUMPED_0;
  wire       [38:0]   decode_ctrls_0_up_Prediction_WORD_JUMP_PC_0;
  wire       [1:0]    decode_ctrls_0_up_Prediction_WORD_SLICES_TAKEN_0;
  wire       [1:0]    decode_ctrls_0_up_Prediction_WORD_SLICES_BRANCH_0;
  wire       [11:0]   decode_ctrls_0_up_Prediction_BRANCH_HISTORY_0;
  wire       [1:0]    decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_0_0;
  wire       [1:0]    decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_0_1;
  wire       [9:0]    decode_ctrls_0_up_Fetch_ID_0;
  wire       [9:0]    decode_ctrls_0_up_Decode_DOP_ID_0;
  wire       [38:0]   decode_ctrls_0_up_PC_0;
  wire       [0:0]    decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0;
  reg        [31:0]   decode_ctrls_0_up_Decode_INSTRUCTION_RAW_0;
  reg                 decode_ctrls_0_up_Decode_DECOMPRESSION_FAULT_0;
  reg        [31:0]   decode_ctrls_0_up_Decode_INSTRUCTION_0;
  wire                decode_ctrls_0_up_isFiring;
  wire       [1:0]    fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_LAST;
  wire                fetch_logic_ctrls_2_down_Prediction_WORD_JUMPED;
  wire       [0:0]    fetch_logic_ctrls_2_down_Prediction_WORD_JUMP_SLICE;
  wire       [1:0]    fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK;
  (* keep , syn_keep *) wire       [38:0]   execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [38:0]   execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) reg        [38:0]   execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0 /* synthesis syn_keep = 1 */ ;
  wire       [0:0]    execute_ctrl2_down_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  wire       [1:0]    execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0;
  wire       [1:0]    execute_ctrl3_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
  wire                execute_ctrl3_down_lane0_IntFormatPlugin_logic_SIGNED_lane0;
  wire       [1:0]    execute_ctrl4_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
  wire                execute_ctrl4_down_lane0_IntFormatPlugin_logic_SIGNED_lane0;
  wire       [1:0]    execute_ctrl2_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
  wire                execute_ctrl2_down_lane0_IntFormatPlugin_logic_SIGNED_lane0;
  wire                execute_ctrl2_down_SrcStageables_UNSIGNED_lane0;
  wire                execute_ctrl2_down_SrcStageables_ZERO_lane0;
  wire                execute_ctrl2_down_SrcStageables_REVERT_lane0;
  wire       [38:0]   execute_ctrl1_down_PC_lane0;
  wire       [63:0]   execute_ctrl1_down_integer_RS2_lane0;
  wire       [1:0]    execute_ctrl1_down_early0_SrcPlugin_logic_SRC2_CTRL_lane0;
  wire       [63:0]   execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0;
  wire       [63:0]   execute_ctrl1_down_integer_RS1_lane0;
  wire       [0:0]    execute_ctrl1_down_early0_SrcPlugin_logic_SRC1_CTRL_lane0;
  wire       [63:0]   execute_ctrl1_down_early0_SrcPlugin_SRC1_lane0;
  wire       [31:0]   execute_ctrl1_down_Decode_UOP_lane0;
  wire                execute_ctrl4_down_AguPlugin_FLOAT_lane0;
  wire       [38:0]   execute_ctrl4_down_PC_lane0;
  wire                execute_ctrl4_down_isReady;
  wire                execute_ctrl4_down_LANE_SEL_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_FROM_ACCESS_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_MMU_FAILURE_lane0;
  reg                 execute_ctrl4_up_COMMIT_lane0;
  wire                execute_ctrl4_down_COMMIT_lane0;
  reg                 execute_ctrl4_COMMIT_lane0_bypass;
  reg                 execute_ctrl4_up_TRAP_lane0;
  wire                execute_ctrl4_down_TRAP_lane0;
  reg                 execute_ctrl4_TRAP_lane0_bypass;
  wire                execute_ctrl4_down_AguPlugin_SEL_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_FROM_PREFETCH_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_FENCE_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_onTrigger_HIT_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0;
  wire                execute_ctrl4_down_MMU_BYPASS_TRANSLATION_lane0;
  wire                execute_ctrl4_down_AguPlugin_STORE_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0;
  wire                execute_ctrl4_down_MMU_HAZARD_lane0;
  wire                execute_ctrl4_down_MMU_REFILL_lane0;
  wire                execute_ctrl4_down_MMU_ACCESS_FAULT_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_MMU_PAGE_FAULT_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_onPma_IO_RSP_lane0_fault;
  wire                execute_ctrl4_down_LsuPlugin_logic_onPma_IO_RSP_lane0_io;
  wire                execute_ctrl4_down_LsuPlugin_logic_pmpPort_ACCESS_FAULT_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault;
  wire                execute_ctrl4_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_io;
  wire                execute_ctrl4_down_LsuPlugin_logic_preCtrl_IS_AMO_lane0;
  wire       [31:0]   execute_ctrl4_down_Decode_UOP_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_onCtrl_SC_MISS_lane0;
  wire       [63:0]   execute_ctrl4_down_LsuPlugin_logic_onCtrl_loadData_RESULT_lane0;
  wire       [15:0]   execute_ctrl4_down_Decode_UOP_ID_lane0;
  wire       [1:0]    execute_ctrl4_down_LsuL1_SIZE_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_onPma_IO_lane0;
  reg        [63:0]   execute_ctrl4_up_integer_RS2_lane0;
  reg                 execute_ctrl3_down_MMU_HAZARD_lane0;
  reg                 execute_ctrl3_down_MMU_REFILL_lane0;
  reg                 execute_ctrl3_down_MMU_ACCESS_FAULT_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_MMU_FAILURE_lane0;
  reg                 execute_ctrl3_down_MMU_ALLOW_READ_lane0;
  reg                 execute_ctrl3_down_MMU_ALLOW_WRITE_lane0;
  wire                execute_ctrl3_down_AguPlugin_STORE_lane0;
  reg                 execute_ctrl3_down_MMU_PAGE_FAULT_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_MMU_PAGE_FAULT_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0;
  wire       [63:0]   execute_ctrl3_down_early0_SrcPlugin_ADD_SUB_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_onPma_IO_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_FROM_PREFETCH_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_FENCE_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_FROM_ACCESS_lane0;
  reg                 execute_ctrl3_down_LsuPlugin_logic_onPma_IO_RSP_lane0_fault;
  wire                execute_ctrl3_down_LsuPlugin_logic_onPma_IO_RSP_lane0_io;
  wire                execute_ctrl3_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault;
  wire                execute_ctrl3_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_io;
  wire                execute_ctrl3_down_LsuPlugin_logic_preCtrl_IS_AMO_lane0;
  wire                execute_ctrl3_down_LsuL1_ATOMIC_lane0;
  wire                execute_ctrl3_down_AguPlugin_SEL_lane0;
  wire                execute_ctrl3_down_LsuL1_INVALID_lane0;
  wire                execute_ctrl3_down_LsuL1_CLEAN_lane0;
  reg                 execute_ctrl3_down_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0;
  reg                 execute_ctrl4_LsuL1_SEL_lane0_bypass;
  wire                execute_ctrl4_down_LsuPlugin_logic_FROM_LSU_lane0;
  reg                 execute_ctrl4_up_LsuL1_SEL_lane0;
  reg                 execute_ctrl3_LsuL1_SEL_lane0_bypass;
  reg                 execute_ctrl3_up_LANE_SEL_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_FROM_LSU_lane0;
  reg                 execute_ctrl3_up_LsuL1_SEL_lane0;
  reg        [31:0]   execute_ctrl3_down_MMU_TRANSLATED_lane0;
  reg                 execute_ctrl2_up_LsuPlugin_logic_FENCE_lane0;
  wire                execute_ctrl2_down_LsuPlugin_logic_FENCE_lane0;
  reg                 execute_ctrl2_LsuPlugin_logic_FENCE_lane0_bypass;
  wire                execute_ctrl2_down_LsuPlugin_logic_FROM_PREFETCH_lane0;
  wire                execute_ctrl2_down_LsuPlugin_logic_FROM_LSU_lane0;
  wire       [11:0]   execute_ctrl2_down_Decode_STORE_ID_lane0;
  wire                execute_ctrl2_down_LsuL1_FLUSH_lane0;
  wire                execute_ctrl2_down_LsuL1_PREFETCH_lane0;
  wire                execute_ctrl2_down_LsuL1_INVALID_lane0;
  wire                execute_ctrl2_down_LsuL1_CLEAN_lane0;
  wire                execute_ctrl2_down_LsuL1_STORE_lane0;
  wire                execute_ctrl2_down_LsuL1_ATOMIC_lane0;
  wire                execute_ctrl2_down_LsuL1_LOAD_lane0;
  wire       [1:0]    execute_ctrl2_down_LsuL1_SIZE_lane0;
  wire       [7:0]    execute_ctrl2_down_LsuL1_MASK_lane0;
  wire                execute_ctrl2_down_LsuL1_SEL_lane0;
  wire                execute_ctrl2_down_AguPlugin_INVALIDATE_lane0;
  wire                execute_ctrl2_down_AguPlugin_CLEAN_lane0;
  wire                execute_ctrl2_down_AguPlugin_ATOMIC_lane0;
  wire                execute_ctrl2_down_AguPlugin_STORE_lane0;
  wire                execute_ctrl2_down_AguPlugin_LOAD_lane0;
  wire       [1:0]    execute_ctrl2_down_AguPlugin_SIZE_lane0;
  wire                execute_ctrl2_down_AguPlugin_SEL_lane0;
  wire       [31:0]   execute_ctrl2_down_Decode_UOP_lane0;
  wire                execute_ctrl2_down_LsuPlugin_logic_FROM_WB_lane0;
  wire                execute_ctrl2_down_LsuPlugin_logic_FROM_ACCESS_lane0;
  wire                execute_ctrl2_down_LsuPlugin_logic_FORCE_PHYSICAL_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_onTrigger_HIT_lane0;
  wire       [1:0]    execute_ctrl3_down_LsuL1_SIZE_lane0;
  wire                execute_ctrl3_down_LsuL1_STORE_lane0;
  wire                execute_ctrl3_down_LsuL1_LOAD_lane0;
  wire                execute_ctrl3_down_LsuL1_FLUSH_lane0;
  wire                execute_ctrl3_down_LsuL1_SEL_lane0;
  wire       [31:0]   execute_ctrl0_down_Decode_UOP_lane0;
  wire       [1:0]    execute_ctrl0_down_AguPlugin_SIZE_lane0;
  wire       [2:0]    execute_ctrl2_down_early0_EnvPlugin_OP_lane0;
  wire       [38:0]   execute_ctrl2_down_PC_lane0;
  wire       [15:0]   execute_ctrl2_down_Decode_UOP_ID_lane0;
  wire                decode_ctrls_1_lane0_upIsCancel;
  wire                decode_ctrls_1_lane0_downIsCancel;
  wire       [9:0]    decode_ctrls_0_down_Decode_DOP_ID_0;
  wire       [9:0]    decode_ctrls_0_down_Fetch_ID_0;
  wire       [38:0]   decode_ctrls_0_down_PC_0;
  wire                decode_ctrls_0_up_isReady;
  wire                decode_ctrls_0_up_LANE_SEL_0;
  wire                decode_ctrls_0_lane0_upIsCancel;
  wire                decode_ctrls_0_lane0_downIsCancel;
  wire       [9:0]    fetch_logic_ctrls_0_down_Fetch_ID;
  reg                 _zz_3;
  reg        [1:0]    BtbPlugin_logic_ras_ptr_pop_aheadValue;
  wire                fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_valid;
  wire       [12:0]   fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_address;
  wire       [1:0]    fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_data_0;
  wire       [1:0]    fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_data_1;
  wire       [12:0]   fetch_logic_ctrls_1_down_GSharePlugin_logic_HASH;
  (* keep , syn_keep *) reg        [1:0]    fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) reg        [1:0]    fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_1 /* synthesis syn_keep = 1 */ ;
  wire                fetch_logic_ctrls_0_down_isReady;
  wire                fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_valid;
  wire       [12:0]   fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_address;
  wire       [1:0]    fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_data_0;
  wire       [1:0]    fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_data_1;
  wire       [11:0]   fetch_logic_ctrls_0_down_Prediction_BRANCH_HISTORY;
  wire       [12:0]   fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH;
  reg                 _zz_4;
  wire                fetch_logic_ctrls_2_up_isMoving;
  wire                fetch_logic_ctrls_2_up_isCanceling;
  wire                fetch_logic_ctrls_2_down_isReady;
  wire                fetch_logic_ctrls_2_down_TRAP;
  wire                fetch_logic_ctrls_2_down_MMU_BYPASS_TRANSLATION;
  wire                fetch_logic_ctrls_2_down_Fetch_PC_FAULT;
  wire                fetch_logic_ctrls_2_down_MMU_HAZARD;
  wire                fetch_logic_ctrls_2_down_MMU_REFILL;
  wire                fetch_logic_ctrls_2_down_MMU_ACCESS_FAULT;
  wire                fetch_logic_ctrls_2_down_MMU_ALLOW_EXECUTE;
  wire                fetch_logic_ctrls_2_down_MMU_PAGE_FAULT;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_ACCESS_FAULT;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HIT;
  wire                fetch_logic_ctrls_2_up_isCancel;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_HAZARD;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_0_loaded;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_0_error;
  wire       [19:0]   fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_0_address;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_1_loaded;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_1_error;
  wire       [19:0]   fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_1_address;
  wire       [38:0]   fetch_logic_ctrls_2_down_Fetch_WORD_PC;
  wire                fetch_logic_ctrls_2_up_isReady;
  wire                fetch_logic_ctrls_2_up_isValid;
  wire       [0:0]    fetch_logic_ctrls_2_down_FetchL1Plugin_logic_PLRU_BYPASSED_0;
  wire       [31:0]   fetch_logic_ctrls_2_down_MMU_TRANSLATED;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HIT;
  wire                fetch_logic_ctrls_1_down_MMU_BYPASS_TRANSLATION;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HITS_0;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HITS_1;
  wire       [2:0]    fetch_logic_ctrls_1_down_MMU_WAYS_OH;
  wire       [31:0]   fetch_logic_ctrls_1_down_MMU_WAYS_PHYSICAL_0;
  wire       [31:0]   fetch_logic_ctrls_1_down_MMU_WAYS_PHYSICAL_1;
  wire       [31:0]   fetch_logic_ctrls_1_down_MMU_WAYS_PHYSICAL_2;
  wire       [5:0]    fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE_ADDRESS;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_HAZARD;
  wire       [31:0]   fetch_logic_ctrls_2_down_FetchL1Plugin_logic_BANKS_MUXES_0;
  wire       [31:0]   fetch_logic_ctrls_2_down_FetchL1Plugin_logic_BANKS_MUXES_1;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_0;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_1;
  wire       [31:0]   fetch_logic_ctrls_2_down_Fetch_WORD;
  wire       [38:0]   fetch_logic_ctrls_1_down_Fetch_WORD_PC;
  wire       [31:0]   fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_0;
  wire       [31:0]   fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_1;
  wire       [0:0]    fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_0;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_VALID;
  reg        [0:0]    fetch_logic_ctrls_1_down_FetchL1Plugin_logic_PLRU_BYPASSED_0;
  wire       [5:0]    fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE_ADDRESS;
  wire                fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE;
  wire       [0:0]    fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_0;
  wire                fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_VALID;
  reg                 fetch_logic_ctrls_1_up_valid;
  wire                fetch_logic_ctrls_1_up_ready;
  wire       [38:0]   fetch_logic_ctrls_0_down_Fetch_WORD_PC;
  reg                 _zz_fetch_logic_ctrls_0_haltRequest_FetchL1Plugin_l217;
  wire       [0:0]    fetch_logic_ctrls_1_down_FetchL1Plugin_logic_PLRU_READ_0;
  reg                 _zz_5;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_loaded;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_error;
  wire       [19:0]   fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_address;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_loaded;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_error;
  wire       [19:0]   fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_address;
  reg                 _zz_6;
  wire       [63:0]   fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_WORDS_0;
  wire       [63:0]   fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_WORDS_1;
  reg                 _zz_7;
  wire                fetch_logic_ctrls_0_down_isFiring;
  wire       [63:0]   execute_ctrl3_down_DivPlugin_DIV_RESULT_lane0;
  wire                execute_ctrl3_down_early0_DivPlugin_SEL_lane0;
  wire       [63:0]   execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0;
  wire                execute_ctrl2_down_early0_DivPlugin_SEL_lane0;
  reg                 execute_ctrl2_up_LANE_SEL_lane0;
  wire                execute_ctrl2_down_isReady;
  wire                execute_ctrl2_down_DivPlugin_REM_lane0;
  wire       [63:0]   execute_ctrl2_down_RsUnsignedPlugin_RS2_UNSIGNED_lane0;
  wire       [63:0]   execute_ctrl2_down_RsUnsignedPlugin_RS1_UNSIGNED_lane0;
  wire                execute_ctrl2_down_RsUnsignedPlugin_RS2_REVERT_lane0;
  wire                execute_ctrl2_down_RsUnsignedPlugin_RS1_REVERT_lane0;
  wire                execute_ctrl2_down_RsUnsignedPlugin_IS_W_lane0;
  reg        [63:0]   execute_ctrl2_down_RsUnsignedPlugin_RS2_FORMATED_lane0;
  reg        [63:0]   execute_ctrl2_down_RsUnsignedPlugin_RS1_FORMATED_lane0;
  wire                execute_ctrl4_down_early0_MulPlugin_SEL_lane0;
  wire                execute_ctrl4_down_MulPlugin_HIGH_lane0;
  wire       [130:0]  execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0;
  wire       [25:0]   execute_ctrl4_down_early0_MulPlugin_logic_steps_0_adders_2_lane0;
  wire       [46:0]   execute_ctrl4_down_early0_MulPlugin_logic_steps_0_adders_1_lane0;
  wire       [63:0]   execute_ctrl4_down_early0_MulPlugin_logic_steps_0_adders_0_lane0;
  wire       [25:0]   execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_15_lane0;
  wire       [42:0]   execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_14_lane0;
  wire       [42:0]   execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_13_lane0;
  wire       [33:0]   execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_12_lane0;
  wire       [59:0]   execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_11_lane0;
  wire       [59:0]   execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_10_lane0;
  wire       [33:0]   execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_9_lane0;
  wire       [33:0]   execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_8_lane0;
  wire       [76:0]   execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_7_lane0;
  wire       [76:0]   execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_6_lane0;
  wire       [33:0]   execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_5_lane0;
  wire       [33:0]   execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_4_lane0;
  wire       [33:0]   execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_3_lane0;
  wire       [33:0]   execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_2_lane0;
  wire       [33:0]   execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_1_lane0;
  wire       [33:0]   execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_0_lane0;
  wire       [25:0]   execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0;
  wire       [46:0]   execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0;
  wire       [63:0]   execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0;
  wire       [25:0]   execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_15_lane0;
  wire       [42:0]   execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_14_lane0;
  wire       [42:0]   execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_13_lane0;
  wire       [33:0]   execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_12_lane0;
  wire       [59:0]   execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_11_lane0;
  wire       [59:0]   execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_10_lane0;
  wire       [33:0]   execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_9_lane0;
  wire       [33:0]   execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_8_lane0;
  wire       [76:0]   execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_7_lane0;
  wire       [76:0]   execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_6_lane0;
  wire       [33:0]   execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_5_lane0;
  wire       [33:0]   execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_4_lane0;
  wire       [33:0]   execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_3_lane0;
  wire       [33:0]   execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_2_lane0;
  wire       [33:0]   execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_1_lane0;
  wire       [33:0]   execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_0_lane0;
  wire       [25:0]   execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_15_lane0;
  wire       [42:0]   execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_14_lane0;
  wire       [42:0]   execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_13_lane0;
  wire       [33:0]   execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_12_lane0;
  wire       [59:0]   execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_11_lane0;
  wire       [59:0]   execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_10_lane0;
  wire       [33:0]   execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_9_lane0;
  wire       [33:0]   execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_8_lane0;
  wire       [76:0]   execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_7_lane0;
  wire       [76:0]   execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_6_lane0;
  wire       [33:0]   execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_5_lane0;
  wire       [33:0]   execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_4_lane0;
  wire       [33:0]   execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_3_lane0;
  wire       [33:0]   execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_2_lane0;
  wire       [33:0]   execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_1_lane0;
  wire       [33:0]   execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_0_lane0;
  wire                execute_ctrl2_down_RsUnsignedPlugin_RS2_SIGNED_lane0;
  wire       [64:0]   execute_ctrl2_down_MUL_SRC2_lane0;
  wire                execute_ctrl2_down_RsUnsignedPlugin_RS1_SIGNED_lane0;
  wire       [64:0]   execute_ctrl2_down_MUL_SRC1_lane0;
  reg        [63:0]   execute_ctrl2_up_integer_RS2_lane0;
  reg        [63:0]   execute_ctrl2_up_integer_RS1_lane0;
  wire       [63:0]   execute_ctrl4_down_LsuL1_READ_DATA_lane0;
  wire       [63:0]   execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0;
  wire       [7:0]    execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0;
  wire       [63:0]   execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0;
  wire       [7:0]    execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0;
  wire       [1:0]    execute_ctrl4_down_LsuL1Plugin_logic_WRITE_TO_READ_HAZARDS_lane0;
  reg        [63:0]   execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0;
  wire       [7:0]    execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0;
  wire       [63:0]   execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0;
  wire                execute_ctrl4_down_LsuL1_FLUSH_HIT_lane0;
  wire                execute_ctrl4_down_LsuL1_CBM_REDO_lane0;
  wire       [7:0]    execute_ctrl4_down_LsuL1_MASK_lane0;
  wire       [63:0]   execute_ctrl4_down_LsuL1_WRITE_DATA_lane0;
  wire       [38:0]   execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0;
  wire       [0:0]    execute_ctrl4_down_LsuL1_WAIT_WRITEBACK_lane0;
  wire       [0:0]    execute_ctrl4_down_LsuL1_WAIT_REFILL_lane0;
  wire                execute_ctrl4_down_LsuL1_SKIP_WRITE_lane0;
  wire                execute_ctrl4_down_LsuL1_INVALID_lane0;
  wire                execute_ctrl4_down_LsuL1_CLEAN_lane0;
  wire                execute_ctrl4_down_LsuL1_SEL_lane0;
  wire                execute_ctrl4_up_isReady;
  reg                 execute_ctrl4_up_LANE_SEL_lane0;
  wire                execute_ctrl4_down_LsuL1_REFILL_HIT_lane0;
  wire                execute_ctrl4_down_LsuL1_MISS_UNIQUE_lane0;
  wire                execute_ctrl4_down_LsuL1_FAULT_lane0;
  wire                execute_ctrl4_down_LsuL1_MISS_lane0;
  wire                execute_ctrl4_down_LsuL1_FLUSH_HAZARD_lane0;
  wire                execute_ctrl4_down_LsuL1_HAZARD_lane0;
  wire                execute_ctrl4_down_LsuL1Plugin_logic_HAZARD_FORCED_lane0;
  wire                execute_ctrl4_down_LsuL1_FLUSH_lane0;
  wire                execute_ctrl4_down_LsuL1_ABORD_lane0;
  wire                execute_ctrl4_down_LsuL1_PREFETCH_lane0;
  wire                execute_ctrl4_down_LsuL1_LOAD_lane0;
  wire       [1:0]    execute_ctrl4_down_LsuL1Plugin_logic_BANK_BUSY_REMAPPED_lane0;
  wire       [31:0]   execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0;
  wire                execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_loaded;
  wire       [19:0]   execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_address;
  wire                execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault;
  wire                execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_loaded;
  wire       [19:0]   execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_address;
  wire                execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault;
  wire       [0:0]    execute_ctrl4_down_LsuL1Plugin_logic_SHARED_lane0_plru_0;
  wire       [1:0]    execute_ctrl4_down_LsuL1Plugin_logic_SHARED_lane0_dirty;
  wire                execute_ctrl4_down_LsuL1_ATOMIC_lane0;
  wire                execute_ctrl4_down_LsuL1_STORE_lane0;
  wire                execute_ctrl4_down_LsuL1Plugin_logic_NEED_UNIQUE_lane0;
  wire                execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HIT_lane0;
  reg        [1:0]    execute_ctrl3_down_LsuL1Plugin_logic_WAYS_HITS_lane0;
  wire       [0:0]    execute_ctrl3_down_LsuL1Plugin_logic_SHARED_lane0_plru_0;
  wire       [1:0]    execute_ctrl3_down_LsuL1Plugin_logic_SHARED_lane0_dirty;
  wire       [0:0]    execute_ctrl3_LsuL1Plugin_logic_SHARED_lane0_bypass_plru_0;
  wire       [1:0]    execute_ctrl3_LsuL1Plugin_logic_SHARED_lane0_bypass_dirty;
  wire       [0:0]    execute_ctrl3_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_plru_0;
  wire       [1:0]    execute_ctrl3_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_dirty;
  wire                execute_ctrl3_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALID_lane0;
  wire                execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_loaded;
  wire       [19:0]   execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_address;
  wire                execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault;
  wire                execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_loaded;
  wire       [19:0]   execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_address;
  wire                execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault;
  reg        [0:0]    execute_ctrl3_up_LsuL1Plugin_logic_SHARED_lane0_plru_0;
  reg        [1:0]    execute_ctrl3_up_LsuL1Plugin_logic_SHARED_lane0_dirty;
  wire       [0:0]    execute_ctrl2_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_plru_0;
  wire       [1:0]    execute_ctrl2_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_dirty;
  wire                execute_ctrl2_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALID_lane0;
  reg                 execute_ctrl4_up_LsuL1Plugin_logic_FREEZE_HAZARD_lane0;
  wire                execute_ctrl4_down_LsuL1Plugin_logic_FREEZE_HAZARD_lane0;
  wire                execute_ctrl4_LsuL1Plugin_logic_FREEZE_HAZARD_lane0_bypass;
  reg                 execute_ctrl3_up_LsuL1Plugin_logic_FREEZE_HAZARD_lane0;
  wire                execute_ctrl3_down_LsuL1Plugin_logic_FREEZE_HAZARD_lane0;
  wire                execute_ctrl3_LsuL1Plugin_logic_FREEZE_HAZARD_lane0_bypass;
  wire                execute_ctrl2_up_LsuL1Plugin_logic_FREEZE_HAZARD_lane0;
  wire       [31:0]   execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_ADDRESS_lane0;
  wire                execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_VALID_lane0;
  wire       [31:0]   execute_ctrl3_down_LsuL1_PHYSICAL_ADDRESS_lane0;
  wire       [31:0]   execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_ADDRESS_lane0;
  wire                execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_VALID_lane0;
  reg        [1:0]    execute_ctrl3_down_LsuL1Plugin_logic_WRITE_TO_READ_HAZARDS_lane0;
  wire       [63:0]   execute_ctrl4_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0;
  wire       [63:0]   execute_ctrl4_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1;
  wire       [1:0]    execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0;
  wire       [63:0]   execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0;
  wire       [38:0]   execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0;
  wire       [63:0]   execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0;
  wire       [63:0]   execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1;
  wire       [1:0]    execute_ctrl3_down_LsuL1Plugin_logic_BANK_BUSY_lane0;
  reg        [1:0]    execute_ctrl3_down_LsuL1Plugin_logic_BANK_BUSY_REMAPPED_lane0;
  wire       [63:0]   execute_ctrl3_down_LsuL1Plugin_logic_BANKS_WORDS_lane0_0;
  wire       [63:0]   execute_ctrl3_down_LsuL1Plugin_logic_BANKS_WORDS_lane0_1;
  reg        [1:0]    execute_ctrl2_down_LsuL1Plugin_logic_BANK_BUSY_lane0;
  wire       [38:0]   execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0;
  reg                 _zz_8;
  reg                 _zz_9;
  wire                execute_ctrl2_down_early0_BarrelShifterPlugin_SEL_lane0;
  wire       [63:0]   execute_ctrl2_down_early0_BarrelShifterPlugin_SHIFT_RESULT_lane0;
  wire                execute_ctrl2_down_BarrelShifterPlugin_IS_W_lane0;
  wire                execute_ctrl2_down_BarrelShifterPlugin_IS_W_RIGHT_lane0;
  wire                execute_ctrl2_down_BarrelShifterPlugin_SIGNED_lane0;
  wire                execute_ctrl2_down_BarrelShifterPlugin_LEFT_lane0;
  wire                execute_ctrl2_down_early0_IntAluPlugin_SEL_lane0;
  wire       [63:0]   execute_ctrl2_down_early0_IntAluPlugin_ALU_RESULT_lane0;
  wire                execute_ctrl2_down_early0_IntAluPlugin_ALU_SLTX_lane0;
  wire                execute_ctrl2_down_early0_SrcPlugin_LESS_lane0;
  wire                execute_ctrl2_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0;
  wire       [63:0]   execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0;
  wire       [63:0]   execute_ctrl2_down_early0_SrcPlugin_SRC2_lane0;
  wire       [63:0]   execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0;
  wire       [1:0]    execute_ctrl2_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  wire                early0_BranchPlugin_logic_events_branchMiss;
  wire                early0_BranchPlugin_logic_events_branchCount;
  reg                 MmuPlugin_api_fetchTranslationEnable;
  reg                 MmuPlugin_api_lsuTranslationEnable;
  wire                AlignerPlugin_api_singleFetch;
  wire                AlignerPlugin_api_downMoving;
  wire                AlignerPlugin_api_haltIt;
  reg                 DispatchPlugin_api_haltDispatch;
  wire                execute_freeze_valid;
  wire       [0:0]    execute_lane0_api_hartsInflight;
  wire                execute_lane0_ctrls_2_upIsCancel;
  wire                execute_lane0_ctrls_2_downIsCancel;
  reg                 CsrRamPlugin_api_holdRead;
  reg                 CsrRamPlugin_api_holdWrite;
  reg                 CsrAccessPlugin_bus_decode_exception;
  wire                CsrAccessPlugin_bus_decode_read;
  wire                CsrAccessPlugin_bus_decode_write;
  wire       [11:0]   CsrAccessPlugin_bus_decode_address;
  reg                 CsrAccessPlugin_bus_decode_trap;
  wire                PrivilegedPlugin_api_lsuTriggerBus_load;
  wire                PrivilegedPlugin_api_lsuTriggerBus_store;
  reg                 TrapPlugin_api_harts_0_redo;
  reg                 TrapPlugin_api_harts_0_askWake;
  reg                 TrapPlugin_api_harts_0_rvTrap;
  wire                TrapPlugin_api_harts_0_fsmBusy;
  wire                TrapPlugin_api_harts_0_holdPrivChange;
  reg                 MmuPlugin_logic_accessBus_cmd_valid;
  wire                MmuPlugin_logic_accessBus_cmd_ready;
  wire       [31:0]   MmuPlugin_logic_accessBus_cmd_payload_address;
  wire       [1:0]    MmuPlugin_logic_accessBus_cmd_payload_size;
  wire                MmuPlugin_logic_accessBus_rsp_valid;
  wire       [63:0]   MmuPlugin_logic_accessBus_rsp_payload_data;
  reg                 MmuPlugin_logic_accessBus_rsp_payload_error;
  reg                 MmuPlugin_logic_accessBus_rsp_payload_redo;
  wire                MmuPlugin_logic_accessBus_rsp_payload_waitAny;
  reg        [3:0]    MmuPlugin_logic_satp_mode;
  reg        [43:0]   MmuPlugin_logic_satp_ppn;
  reg                 MmuPlugin_logic_status_mxr;
  reg                 MmuPlugin_logic_status_sum;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_1;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_2;
  wire                PmpPlugin_logic_entries_0_isLocked;
  reg        [20:0]   PmpPlugin_logic_entries_0_address;
  reg        [1:0]    PmpPlugin_logic_entries_0_cfg_kind;
  reg                 PmpPlugin_logic_entries_0_cfg_read;
  reg                 PmpPlugin_logic_entries_0_cfg_write;
  reg                 PmpPlugin_logic_entries_0_cfg_execute;
  reg                 PmpPlugin_logic_entries_0_cfg_locked;
  reg        [1:0]    PmpPlugin_logic_entries_0_cfgNext_kind;
  reg                 PmpPlugin_logic_entries_0_cfgNext_read;
  reg                 PmpPlugin_logic_entries_0_cfgNext_write;
  reg                 PmpPlugin_logic_entries_0_cfgNext_execute;
  reg                 PmpPlugin_logic_entries_0_cfgNext_locked;
  wire                when_PmpPlugin_l127;
  wire                when_PmpPlugin_l129;
  reg                 PmpPlugin_logic_entries_0_isNapot;
  reg                 PmpPlugin_logic_entries_0_isTor;
  wire       [19:0]   _zz_PmpPlugin_logic_entries_0_napot;
  wire                _zz_PmpPlugin_logic_entries_0_napot_1;
  wire                _zz_PmpPlugin_logic_entries_0_napot_2;
  wire                _zz_PmpPlugin_logic_entries_0_napot_3;
  wire                _zz_PmpPlugin_logic_entries_0_napot_4;
  wire                _zz_PmpPlugin_logic_entries_0_napot_5;
  wire                _zz_PmpPlugin_logic_entries_0_napot_6;
  wire                _zz_PmpPlugin_logic_entries_0_napot_7;
  wire                _zz_PmpPlugin_logic_entries_0_napot_8;
  wire                _zz_PmpPlugin_logic_entries_0_napot_9;
  wire                _zz_PmpPlugin_logic_entries_0_napot_10;
  wire                _zz_PmpPlugin_logic_entries_0_napot_11;
  wire                _zz_PmpPlugin_logic_entries_0_napot_12;
  wire                _zz_PmpPlugin_logic_entries_0_napot_13;
  wire                _zz_PmpPlugin_logic_entries_0_napot_14;
  wire                _zz_PmpPlugin_logic_entries_0_napot_15;
  reg        [19:0]   _zz_PmpPlugin_logic_entries_0_napot_16;
  wire                _zz_PmpPlugin_logic_entries_0_napot_17;
  wire                _zz_PmpPlugin_logic_entries_0_napot_18;
  wire                _zz_PmpPlugin_logic_entries_0_napot_19;
  wire                _zz_PmpPlugin_logic_entries_0_napot_20;
  wire                _zz_PmpPlugin_logic_entries_0_napot_21;
  wire                _zz_PmpPlugin_logic_entries_0_napot_22;
  wire                _zz_PmpPlugin_logic_entries_0_napot_23;
  wire       [19:0]   PmpPlugin_logic_entries_0_napot;
  reg        [19:0]   PmpPlugin_logic_entries_0_mask;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3;
  reg        [9:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5;
  wire                PmpPlugin_logic_entries_1_isLocked;
  reg        [20:0]   PmpPlugin_logic_entries_1_address;
  reg        [1:0]    PmpPlugin_logic_entries_1_cfg_kind;
  reg                 PmpPlugin_logic_entries_1_cfg_read;
  reg                 PmpPlugin_logic_entries_1_cfg_write;
  reg                 PmpPlugin_logic_entries_1_cfg_execute;
  reg                 PmpPlugin_logic_entries_1_cfg_locked;
  reg        [1:0]    PmpPlugin_logic_entries_1_cfgNext_kind;
  reg                 PmpPlugin_logic_entries_1_cfgNext_read;
  reg                 PmpPlugin_logic_entries_1_cfgNext_write;
  reg                 PmpPlugin_logic_entries_1_cfgNext_execute;
  reg                 PmpPlugin_logic_entries_1_cfgNext_locked;
  wire                when_PmpPlugin_l127_1;
  wire                when_PmpPlugin_l129_1;
  reg                 PmpPlugin_logic_entries_1_isNapot;
  reg                 PmpPlugin_logic_entries_1_isTor;
  wire       [19:0]   _zz_PmpPlugin_logic_entries_1_napot;
  wire                _zz_PmpPlugin_logic_entries_1_napot_1;
  wire                _zz_PmpPlugin_logic_entries_1_napot_2;
  wire                _zz_PmpPlugin_logic_entries_1_napot_3;
  wire                _zz_PmpPlugin_logic_entries_1_napot_4;
  wire                _zz_PmpPlugin_logic_entries_1_napot_5;
  wire                _zz_PmpPlugin_logic_entries_1_napot_6;
  wire                _zz_PmpPlugin_logic_entries_1_napot_7;
  wire                _zz_PmpPlugin_logic_entries_1_napot_8;
  wire                _zz_PmpPlugin_logic_entries_1_napot_9;
  wire                _zz_PmpPlugin_logic_entries_1_napot_10;
  wire                _zz_PmpPlugin_logic_entries_1_napot_11;
  wire                _zz_PmpPlugin_logic_entries_1_napot_12;
  wire                _zz_PmpPlugin_logic_entries_1_napot_13;
  wire                _zz_PmpPlugin_logic_entries_1_napot_14;
  wire                _zz_PmpPlugin_logic_entries_1_napot_15;
  reg        [19:0]   _zz_PmpPlugin_logic_entries_1_napot_16;
  wire                _zz_PmpPlugin_logic_entries_1_napot_17;
  wire                _zz_PmpPlugin_logic_entries_1_napot_18;
  wire                _zz_PmpPlugin_logic_entries_1_napot_19;
  wire                _zz_PmpPlugin_logic_entries_1_napot_20;
  wire                _zz_PmpPlugin_logic_entries_1_napot_21;
  wire                _zz_PmpPlugin_logic_entries_1_napot_22;
  wire                _zz_PmpPlugin_logic_entries_1_napot_23;
  wire       [19:0]   PmpPlugin_logic_entries_1_napot;
  reg        [19:0]   PmpPlugin_logic_entries_1_mask;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_6;
  reg        [9:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_7;
  wire                PmpPlugin_logic_entries_2_isLocked;
  reg        [20:0]   PmpPlugin_logic_entries_2_address;
  reg        [1:0]    PmpPlugin_logic_entries_2_cfg_kind;
  reg                 PmpPlugin_logic_entries_2_cfg_read;
  reg                 PmpPlugin_logic_entries_2_cfg_write;
  reg                 PmpPlugin_logic_entries_2_cfg_execute;
  reg                 PmpPlugin_logic_entries_2_cfg_locked;
  reg        [1:0]    PmpPlugin_logic_entries_2_cfgNext_kind;
  reg                 PmpPlugin_logic_entries_2_cfgNext_read;
  reg                 PmpPlugin_logic_entries_2_cfgNext_write;
  reg                 PmpPlugin_logic_entries_2_cfgNext_execute;
  reg                 PmpPlugin_logic_entries_2_cfgNext_locked;
  wire                when_PmpPlugin_l127_2;
  wire                when_PmpPlugin_l129_2;
  reg                 PmpPlugin_logic_entries_2_isNapot;
  reg                 PmpPlugin_logic_entries_2_isTor;
  wire       [19:0]   _zz_PmpPlugin_logic_entries_2_napot;
  wire                _zz_PmpPlugin_logic_entries_2_napot_1;
  wire                _zz_PmpPlugin_logic_entries_2_napot_2;
  wire                _zz_PmpPlugin_logic_entries_2_napot_3;
  wire                _zz_PmpPlugin_logic_entries_2_napot_4;
  wire                _zz_PmpPlugin_logic_entries_2_napot_5;
  wire                _zz_PmpPlugin_logic_entries_2_napot_6;
  wire                _zz_PmpPlugin_logic_entries_2_napot_7;
  wire                _zz_PmpPlugin_logic_entries_2_napot_8;
  wire                _zz_PmpPlugin_logic_entries_2_napot_9;
  wire                _zz_PmpPlugin_logic_entries_2_napot_10;
  wire                _zz_PmpPlugin_logic_entries_2_napot_11;
  wire                _zz_PmpPlugin_logic_entries_2_napot_12;
  wire                _zz_PmpPlugin_logic_entries_2_napot_13;
  wire                _zz_PmpPlugin_logic_entries_2_napot_14;
  wire                _zz_PmpPlugin_logic_entries_2_napot_15;
  reg        [19:0]   _zz_PmpPlugin_logic_entries_2_napot_16;
  wire                _zz_PmpPlugin_logic_entries_2_napot_17;
  wire                _zz_PmpPlugin_logic_entries_2_napot_18;
  wire                _zz_PmpPlugin_logic_entries_2_napot_19;
  wire                _zz_PmpPlugin_logic_entries_2_napot_20;
  wire                _zz_PmpPlugin_logic_entries_2_napot_21;
  wire                _zz_PmpPlugin_logic_entries_2_napot_22;
  wire                _zz_PmpPlugin_logic_entries_2_napot_23;
  wire       [19:0]   PmpPlugin_logic_entries_2_napot;
  reg        [19:0]   PmpPlugin_logic_entries_2_mask;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_8;
  reg        [9:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_9;
  wire                PmpPlugin_logic_entries_3_isLocked;
  reg        [20:0]   PmpPlugin_logic_entries_3_address;
  reg        [1:0]    PmpPlugin_logic_entries_3_cfg_kind;
  reg                 PmpPlugin_logic_entries_3_cfg_read;
  reg                 PmpPlugin_logic_entries_3_cfg_write;
  reg                 PmpPlugin_logic_entries_3_cfg_execute;
  reg                 PmpPlugin_logic_entries_3_cfg_locked;
  reg        [1:0]    PmpPlugin_logic_entries_3_cfgNext_kind;
  reg                 PmpPlugin_logic_entries_3_cfgNext_read;
  reg                 PmpPlugin_logic_entries_3_cfgNext_write;
  reg                 PmpPlugin_logic_entries_3_cfgNext_execute;
  reg                 PmpPlugin_logic_entries_3_cfgNext_locked;
  wire                when_PmpPlugin_l127_3;
  wire                when_PmpPlugin_l129_3;
  reg                 PmpPlugin_logic_entries_3_isNapot;
  reg                 PmpPlugin_logic_entries_3_isTor;
  wire       [19:0]   _zz_PmpPlugin_logic_entries_3_napot;
  wire                _zz_PmpPlugin_logic_entries_3_napot_1;
  wire                _zz_PmpPlugin_logic_entries_3_napot_2;
  wire                _zz_PmpPlugin_logic_entries_3_napot_3;
  wire                _zz_PmpPlugin_logic_entries_3_napot_4;
  wire                _zz_PmpPlugin_logic_entries_3_napot_5;
  wire                _zz_PmpPlugin_logic_entries_3_napot_6;
  wire                _zz_PmpPlugin_logic_entries_3_napot_7;
  wire                _zz_PmpPlugin_logic_entries_3_napot_8;
  wire                _zz_PmpPlugin_logic_entries_3_napot_9;
  wire                _zz_PmpPlugin_logic_entries_3_napot_10;
  wire                _zz_PmpPlugin_logic_entries_3_napot_11;
  wire                _zz_PmpPlugin_logic_entries_3_napot_12;
  wire                _zz_PmpPlugin_logic_entries_3_napot_13;
  wire                _zz_PmpPlugin_logic_entries_3_napot_14;
  wire                _zz_PmpPlugin_logic_entries_3_napot_15;
  reg        [19:0]   _zz_PmpPlugin_logic_entries_3_napot_16;
  wire                _zz_PmpPlugin_logic_entries_3_napot_17;
  wire                _zz_PmpPlugin_logic_entries_3_napot_18;
  wire                _zz_PmpPlugin_logic_entries_3_napot_19;
  wire                _zz_PmpPlugin_logic_entries_3_napot_20;
  wire                _zz_PmpPlugin_logic_entries_3_napot_21;
  wire                _zz_PmpPlugin_logic_entries_3_napot_22;
  wire                _zz_PmpPlugin_logic_entries_3_napot_23;
  wire       [19:0]   PmpPlugin_logic_entries_3_napot;
  reg        [19:0]   PmpPlugin_logic_entries_3_mask;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_10;
  reg        [9:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_11;
  wire                BtbPlugin_logic_pcPort_valid;
  wire                BtbPlugin_logic_pcPort_payload_fault;
  wire       [38:0]   BtbPlugin_logic_pcPort_payload_pc;
  wire                PcPlugin_logic_harts_0_aggregator_sortedByPriority_2_laneValid;
  wire                BtbPlugin_logic_historyPort_valid;
  wire       [11:0]   BtbPlugin_logic_historyPort_payload_history;
  wire                BtbPlugin_logic_flushPort_valid;
  wire                BtbPlugin_logic_flushPort_payload_self;
  wire                FetchL1Plugin_logic_bus_cmd_valid;
  wire                FetchL1Plugin_logic_bus_cmd_ready;
  wire       [31:0]   FetchL1Plugin_logic_bus_cmd_payload_address;
  wire                FetchL1Plugin_logic_bus_cmd_payload_io;
  wire                FetchL1Plugin_logic_bus_rsp_valid;
  wire                FetchL1Plugin_logic_bus_rsp_ready;
  wire       [63:0]   FetchL1Plugin_logic_bus_rsp_payload_data;
  wire                FetchL1Plugin_logic_bus_rsp_payload_error;
  reg                 FetchL1Plugin_logic_trapPort_valid;
  reg                 FetchL1Plugin_logic_trapPort_payload_exception;
  wire       [38:0]   FetchL1Plugin_logic_trapPort_payload_tval;
  wire       [0:0]    decode_logic_trapPending;
  wire       [0:0]    DispatchPlugin_logic_trapPendings;
  wire       [0:0]    execute_lane0_logic_trapPending;
  wire                early0_IntAluPlugin_logic_wb_valid;
  wire       [63:0]   early0_IntAluPlugin_logic_wb_payload;
  (* keep , syn_keep *) reg        [63:0]   early0_IntAluPlugin_logic_alu_bitwise /* synthesis syn_keep = 1 */ ;
  wire       [63:0]   early0_IntAluPlugin_logic_alu_result;
  wire                early0_BarrelShifterPlugin_logic_wb_valid;
  wire       [63:0]   early0_BarrelShifterPlugin_logic_wb_payload;
  reg        [5:0]    early0_BarrelShifterPlugin_logic_shift_amplitude;
  reg        [63:0]   early0_BarrelShifterPlugin_logic_shift_reversed;
  wire       [63:0]   early0_BarrelShifterPlugin_logic_shift_shifted;
  wire       [63:0]   early0_BarrelShifterPlugin_logic_shift_patched;
  wire                early0_BranchPlugin_logic_wb_valid;
  wire       [63:0]   early0_BranchPlugin_logic_wb_payload;
  wire                early0_BranchPlugin_logic_pcPort_valid;
  wire                early0_BranchPlugin_logic_pcPort_payload_fault;
  wire       [38:0]   early0_BranchPlugin_logic_pcPort_payload_pc;
  wire                PcPlugin_logic_harts_0_aggregator_sortedByPriority_1_laneValid;
  wire                early0_BranchPlugin_logic_historyPort_valid;
  wire       [11:0]   early0_BranchPlugin_logic_historyPort_payload_history;
  wire                early0_BranchPlugin_logic_flushPort_valid;
  reg                 LsuPlugin_logic_events_waiting;
  reg                 LsuPlugin_logic_trapPort_valid;
  reg                 LsuPlugin_logic_trapPort_payload_exception;
  wire       [38:0]   LsuPlugin_logic_trapPort_payload_tval;
  wire                LsuL1_lockPort_valid;
  wire       [31:0]   LsuL1_lockPort_address;
  reg                 LsuL1_ackUnlock;
  wire                LsuL1Plugin_logic_events_loadAccess;
  wire                LsuL1Plugin_logic_events_loadMiss;
  wire                LsuL1Plugin_logic_bus_read_cmd_valid;
  wire                LsuL1Plugin_logic_bus_read_cmd_ready;
  wire       [31:0]   LsuL1Plugin_logic_bus_read_cmd_payload_address;
  wire                LsuL1Plugin_logic_bus_read_rsp_valid;
  wire                LsuL1Plugin_logic_bus_read_rsp_ready;
  wire       [63:0]   LsuL1Plugin_logic_bus_read_rsp_payload_data;
  wire                LsuL1Plugin_logic_bus_read_rsp_payload_error;
  wire                LsuL1Plugin_logic_bus_write_cmd_valid;
  reg                 LsuL1Plugin_logic_bus_write_cmd_ready;
  wire                LsuL1Plugin_logic_bus_write_cmd_payload_last;
  wire       [31:0]   LsuL1Plugin_logic_bus_write_cmd_payload_fragment_address;
  wire       [63:0]   LsuL1Plugin_logic_bus_write_cmd_payload_fragment_data;
  wire                LsuL1Plugin_logic_bus_write_rsp_valid;
  wire                LsuL1Plugin_logic_bus_write_rsp_payload_error;
  reg        [0:0]    LsuL1Plugin_logic_refillCompletions;
  wire                LsuL1Plugin_logic_writebackBusy;
  reg        [1:0]    LsuL1Plugin_logic_banksWrite_mask;
  reg        [8:0]    LsuL1Plugin_logic_banksWrite_address;
  reg        [63:0]   LsuL1Plugin_logic_banksWrite_writeData;
  reg        [7:0]    LsuL1Plugin_logic_banksWrite_writeMask;
  reg        [1:0]    LsuL1Plugin_logic_waysWrite_mask;
  reg        [5:0]    LsuL1Plugin_logic_waysWrite_address;
  reg                 LsuL1Plugin_logic_waysWrite_tag_loaded;
  reg        [19:0]   LsuL1Plugin_logic_waysWrite_tag_address;
  reg                 LsuL1Plugin_logic_waysWrite_tag_fault;
  wire                LsuL1Plugin_logic_waysWrite_valid;
  wire                LsuL1Plugin_logic_banks_0_usedByWriteback;
  wire                LsuL1Plugin_logic_banks_0_write_valid;
  wire       [8:0]    LsuL1Plugin_logic_banks_0_write_payload_address;
  wire       [63:0]   LsuL1Plugin_logic_banks_0_write_payload_data;
  wire       [7:0]    LsuL1Plugin_logic_banks_0_write_payload_mask;
  reg                 LsuL1Plugin_logic_banks_0_read_cmd_valid;
  reg        [8:0]    LsuL1Plugin_logic_banks_0_read_cmd_payload;
  (* keep , syn_keep *) wire       [63:0]   LsuL1Plugin_logic_banks_0_read_rsp /* synthesis syn_keep = 1 */ ;
  wire                LsuL1Plugin_logic_banks_1_usedByWriteback;
  wire                LsuL1Plugin_logic_banks_1_write_valid;
  wire       [8:0]    LsuL1Plugin_logic_banks_1_write_payload_address;
  wire       [63:0]   LsuL1Plugin_logic_banks_1_write_payload_data;
  wire       [7:0]    LsuL1Plugin_logic_banks_1_write_payload_mask;
  reg                 LsuL1Plugin_logic_banks_1_read_cmd_valid;
  reg        [8:0]    LsuL1Plugin_logic_banks_1_read_cmd_payload;
  (* keep , syn_keep *) wire       [63:0]   LsuL1Plugin_logic_banks_1_read_rsp /* synthesis syn_keep = 1 */ ;
  wire                LsuL1Plugin_logic_ways_0_lsuRead_cmd_valid;
  wire       [5:0]    LsuL1Plugin_logic_ways_0_lsuRead_cmd_payload;
  (* keep , syn_keep *) wire                LsuL1Plugin_logic_ways_0_lsuRead_rsp_loaded /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [19:0]   LsuL1Plugin_logic_ways_0_lsuRead_rsp_address /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                LsuL1Plugin_logic_ways_0_lsuRead_rsp_fault /* synthesis syn_keep = 1 */ ;
  wire       [21:0]   _zz_LsuL1Plugin_logic_ways_0_lsuRead_rsp_loaded;
  wire                LsuL1Plugin_logic_ways_1_lsuRead_cmd_valid;
  wire       [5:0]    LsuL1Plugin_logic_ways_1_lsuRead_cmd_payload;
  (* keep , syn_keep *) wire                LsuL1Plugin_logic_ways_1_lsuRead_rsp_loaded /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [19:0]   LsuL1Plugin_logic_ways_1_lsuRead_rsp_address /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                LsuL1Plugin_logic_ways_1_lsuRead_rsp_fault /* synthesis syn_keep = 1 */ ;
  wire       [21:0]   _zz_LsuL1Plugin_logic_ways_1_lsuRead_rsp_loaded;
  reg                 LsuL1Plugin_logic_shared_write_valid;
  reg        [5:0]    LsuL1Plugin_logic_shared_write_payload_address;
  reg        [0:0]    LsuL1Plugin_logic_shared_write_payload_data_plru_0;
  reg        [1:0]    LsuL1Plugin_logic_shared_write_payload_data_dirty;
  wire                LsuL1Plugin_logic_shared_lsuRead_cmd_valid;
  wire       [5:0]    LsuL1Plugin_logic_shared_lsuRead_cmd_payload;
  (* keep , syn_keep *) wire       [0:0]    LsuL1Plugin_logic_shared_lsuRead_rsp_plru_0 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [1:0]    LsuL1Plugin_logic_shared_lsuRead_rsp_dirty /* synthesis syn_keep = 1 */ ;
  wire       [2:0]    _zz_LsuL1Plugin_logic_shared_lsuRead_rsp_plru_0;
  wire                LsuL1Plugin_logic_slotsFreezeHazard;
  wire                LsuL1Plugin_logic_slotsFreeze;
  reg                 LsuL1Plugin_logic_refill_slots_0_valid;
  reg        [31:0]   LsuL1Plugin_logic_refill_slots_0_address;
  reg        [0:0]    LsuL1Plugin_logic_refill_slots_0_way;
  reg                 LsuL1Plugin_logic_refill_slots_0_cmdSent;
  reg                 LsuL1Plugin_logic_refill_slots_0_loadedSet;
  reg                 LsuL1Plugin_logic_refill_slots_0_loaded;
  reg        [0:0]    LsuL1Plugin_logic_refill_slots_0_loadedCounter;
  wire                LsuL1Plugin_logic_refill_slots_0_loadedDone;
  wire                LsuL1Plugin_logic_refill_slots_0_free;
  wire                LsuL1Plugin_logic_refill_slots_0_fire;
  reg        [0:0]    LsuL1Plugin_logic_refill_slots_0_victim;
  wire       [0:0]    LsuL1Plugin_logic_refill_free;
  wire                LsuL1Plugin_logic_refill_full;
  reg                 LsuL1Plugin_logic_refill_push_valid;
  wire       [31:0]   LsuL1Plugin_logic_refill_push_payload_address;
  reg        [0:0]    LsuL1Plugin_logic_refill_push_payload_way;
  reg        [0:0]    LsuL1Plugin_logic_refill_push_payload_victim;
  wire                LsuL1Plugin_logic_refill_push_payload_unique;
  wire                LsuL1Plugin_logic_refill_push_payload_data;
  reg        [31:0]   LsuL1Plugin_logic_refill_pushCounter;
  wire                when_LsuL1Plugin_l382;
  wire                when_LsuL1Plugin_l386;
  wire                LsuL1Plugin_logic_refill_read_arbiter_slotsWithId_0_0;
  wire       [0:0]    LsuL1Plugin_logic_refill_read_arbiter_hits;
  wire                LsuL1Plugin_logic_refill_read_arbiter_hit;
  reg        [0:0]    LsuL1Plugin_logic_refill_read_arbiter_oh;
  reg        [0:0]    LsuL1Plugin_logic_refill_read_arbiter_lock;
  wire                when_LsuL1Plugin_l303;
  wire                LsuL1Plugin_logic_bus_read_cmd_fire;
  wire       [31:0]   LsuL1Plugin_logic_refill_read_cmdAddress;
  wire       [31:0]   LsuL1Plugin_logic_refill_read_rspAddress;
  wire       [0:0]    LsuL1Plugin_logic_refill_read_way;
  (* keep , syn_keep *) reg        [2:0]    LsuL1Plugin_logic_refill_read_wordIndex /* synthesis syn_keep = 1 */ ;
  wire                LsuL1Plugin_logic_refill_read_rspWithData;
  reg        [1:0]    LsuL1Plugin_logic_refill_read_bankWriteNotif;
  wire                LsuL1Plugin_logic_refill_read_writeReservation_win;
  reg                 LsuL1Plugin_logic_refill_read_writeReservation_take;
  reg                 LsuL1Plugin_logic_refill_read_hadError;
  wire                when_LsuL1Plugin_l453;
  reg                 LsuL1Plugin_logic_refill_read_fire;
  wire                LsuL1Plugin_logic_refill_read_reservation_win;
  reg                 LsuL1Plugin_logic_refill_read_reservation_take;
  wire                LsuL1Plugin_logic_refill_read_faulty;
  wire                when_LsuL1Plugin_l466;
  wire       [0:0]    LsuL1_REFILL_BUSY;
  reg                 LsuL1Plugin_logic_writeback_slots_0_fire;
  reg                 LsuL1Plugin_logic_writeback_slots_0_valid;
  reg                 LsuL1Plugin_logic_writeback_slots_0_busy;
  reg        [31:0]   LsuL1Plugin_logic_writeback_slots_0_address;
  reg        [0:0]    LsuL1Plugin_logic_writeback_slots_0_way;
  reg                 LsuL1Plugin_logic_writeback_slots_0_readCmdDone;
  reg                 LsuL1Plugin_logic_writeback_slots_0_readRspDone;
  reg                 LsuL1Plugin_logic_writeback_slots_0_victimBufferReady;
  reg                 LsuL1Plugin_logic_writeback_slots_0_writeCmdDone;
  reg        [0:0]    LsuL1Plugin_logic_writeback_slots_0_timer_counter;
  wire                LsuL1Plugin_logic_writeback_slots_0_timer_done;
  wire                when_LsuL1Plugin_l533;
  wire                LsuL1Plugin_logic_writeback_slots_0_free;
  wire       [0:0]    LsuL1_WRITEBACK_BUSY;
  wire       [0:0]    LsuL1Plugin_logic_writeback_free;
  wire                LsuL1Plugin_logic_writeback_full;
  reg                 LsuL1Plugin_logic_writeback_push_valid;
  reg        [31:0]   LsuL1Plugin_logic_writeback_push_payload_address;
  reg        [0:0]    LsuL1Plugin_logic_writeback_push_payload_way;
  wire                when_LsuL1Plugin_l559;
  wire                when_LsuL1Plugin_l564;
  wire                LsuL1Plugin_logic_writeback_read_arbiter_slotsWithId_0_0;
  wire       [0:0]    LsuL1Plugin_logic_writeback_read_arbiter_hits;
  wire                LsuL1Plugin_logic_writeback_read_arbiter_hit;
  reg        [0:0]    LsuL1Plugin_logic_writeback_read_arbiter_oh;
  reg        [0:0]    LsuL1Plugin_logic_writeback_read_arbiter_lock;
  wire                when_LsuL1Plugin_l303_1;
  wire       [31:0]   LsuL1Plugin_logic_writeback_read_address;
  wire       [0:0]    LsuL1Plugin_logic_writeback_read_way;
  (* keep , syn_keep *) reg        [2:0]    LsuL1Plugin_logic_writeback_read_wordIndex /* synthesis syn_keep = 1 */ ;
  wire                LsuL1Plugin_logic_writeback_read_slotRead_valid;
  wire                LsuL1Plugin_logic_writeback_read_slotRead_payload_last;
  wire       [2:0]    LsuL1Plugin_logic_writeback_read_slotRead_payload_wordIndex;
  wire       [0:0]    LsuL1Plugin_logic_writeback_read_slotRead_payload_way;
  wire                when_LsuL1Plugin_l608;
  reg                 LsuL1Plugin_logic_writeback_read_slotReadLast_valid;
  reg                 LsuL1Plugin_logic_writeback_read_slotReadLast_payload_last;
  reg        [2:0]    LsuL1Plugin_logic_writeback_read_slotReadLast_payload_wordIndex;
  reg        [0:0]    LsuL1Plugin_logic_writeback_read_slotReadLast_payload_way;
  wire       [63:0]   LsuL1Plugin_logic_writeback_read_readedData;
  wire                LsuL1Plugin_logic_writeback_write_arbiter_slotsWithId_0_0;
  wire       [0:0]    LsuL1Plugin_logic_writeback_write_arbiter_hits;
  wire                LsuL1Plugin_logic_writeback_write_arbiter_hit;
  reg        [0:0]    LsuL1Plugin_logic_writeback_write_arbiter_oh;
  reg        [0:0]    LsuL1Plugin_logic_writeback_write_arbiter_lock;
  wire                when_LsuL1Plugin_l303_2;
  (* keep , syn_keep *) reg        [2:0]    LsuL1Plugin_logic_writeback_write_wordIndex /* synthesis syn_keep = 1 */ ;
  wire                LsuL1Plugin_logic_writeback_write_last;
  wire                LsuL1Plugin_logic_writeback_write_bufferRead_valid;
  reg                 LsuL1Plugin_logic_writeback_write_bufferRead_ready;
  wire       [31:0]   LsuL1Plugin_logic_writeback_write_bufferRead_payload_address;
  wire                LsuL1Plugin_logic_writeback_write_bufferRead_payload_last;
  wire                LsuL1Plugin_logic_writeback_write_bufferRead_fire;
  wire                when_LsuL1Plugin_l679;
  wire                LsuL1Plugin_logic_writeback_write_cmd_valid;
  wire                LsuL1Plugin_logic_writeback_write_cmd_ready;
  wire       [31:0]   LsuL1Plugin_logic_writeback_write_cmd_payload_address;
  wire                LsuL1Plugin_logic_writeback_write_cmd_payload_last;
  reg                 LsuL1Plugin_logic_writeback_write_bufferRead_rValid;
  reg        [31:0]   LsuL1Plugin_logic_writeback_write_bufferRead_rData_address;
  reg                 LsuL1Plugin_logic_writeback_write_bufferRead_rData_last;
  wire                when_Stream_l477;
  wire       [2:0]    _zz_LsuL1Plugin_logic_writeback_write_word;
  wire       [63:0]   LsuL1Plugin_logic_writeback_write_word;
  wire       [8:0]    LsuL1Plugin_logic_lsu_rb0_readAddress;
  wire                when_LsuL1Plugin_l721;
  wire                when_LsuL1Plugin_l722;
  wire                when_LsuL1Plugin_l721_1;
  wire                when_LsuL1Plugin_l722_1;
  wire                execute_lane0_ctrls_3_upIsCancel;
  wire                execute_lane0_ctrls_3_downIsCancel;
  reg                 LsuL1Plugin_logic_lsu_rb1_onBanks_0_busyReg;
  wire                when_LsuL1Plugin_l738;
  reg                 LsuL1Plugin_logic_lsu_rb1_onBanks_1_busyReg;
  wire                when_LsuL1Plugin_l738_1;
  wire                execute_lane0_ctrls_4_upIsCancel;
  wire                execute_lane0_ctrls_4_downIsCancel;
  wire                _zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0;
  wire                _zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0_1;
  wire                LsuL1Plugin_logic_lsu_sharedBypassers_0_hit;
  wire       [0:0]    LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_context_state_0;
  wire       [0:0]    LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_evict_id;
  reg        [0:0]    LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_update_id;
  wire       [0:0]    LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_update_state_0;
  wire                LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_evict_sel_0;
  wire                LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_evict_logic_0_state;
  wire                LsuL1Plugin_logic_lsu_ctrl_wayWriteReservation_win;
  reg                 LsuL1Plugin_logic_lsu_ctrl_wayWriteReservation_take;
  wire                LsuL1Plugin_logic_lsu_ctrl_bankWriteReservation_win;
  wire                LsuL1Plugin_logic_lsu_ctrl_bankWriteReservation_take;
  wire       [0:0]    LsuL1Plugin_logic_lsu_ctrl_refillWayWithoutUpdate;
  wire                LsuL1Plugin_logic_lsu_ctrl_refillWayNeedWriteback;
  wire       [0:0]    LsuL1Plugin_logic_lsu_ctrl_refillHazards;
  wire       [0:0]    LsuL1Plugin_logic_lsu_ctrl_writebackHazards;
  wire                LsuL1Plugin_logic_lsu_ctrl_refillHazard;
  wire                LsuL1Plugin_logic_lsu_ctrl_writebackHazard;
  wire                LsuL1Plugin_logic_lsu_ctrl_wasDirty;
  wire       [1:0]    LsuL1Plugin_logic_lsu_ctrl_loadedDirties;
  wire                LsuL1Plugin_logic_lsu_ctrl_refillWayWasDirty;
  wire                LsuL1Plugin_logic_lsu_ctrl_writeToReadHazard;
  wire                LsuL1Plugin_logic_lsu_ctrl_bankNotRead;
  wire                LsuL1Plugin_logic_lsu_ctrl_loadHazard;
  wire                LsuL1Plugin_logic_lsu_ctrl_storeHazard;
  wire                LsuL1Plugin_logic_lsu_ctrl_preventSideEffects;
  wire                LsuL1Plugin_logic_lsu_ctrl_flushHazard;
  wire                LsuL1Plugin_logic_lsu_ctrl_coherencyHazard;
  reg                 LsuL1Plugin_logic_lsu_ctrl_hazardReg;
  reg                 LsuL1Plugin_logic_lsu_ctrl_flushHazardReg;
  wire                LsuL1Plugin_logic_lsu_ctrl_canRefill;
  wire                LsuL1Plugin_logic_lsu_ctrl_canFlush;
  wire       [1:0]    LsuL1Plugin_logic_lsu_ctrl_needFlushs;
  wire       [1:0]    _zz_LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_0;
  wire                LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_0;
  wire                LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_1;
  reg        [1:0]    _zz_LsuL1Plugin_logic_lsu_ctrl_needFlushOh;
  wire       [1:0]    LsuL1Plugin_logic_lsu_ctrl_needFlushOh;
  wire                _zz_LsuL1Plugin_logic_lsu_ctrl_needFlushSel;
  wire       [0:0]    LsuL1Plugin_logic_lsu_ctrl_needFlushSel;
  wire                LsuL1Plugin_logic_lsu_ctrl_isAccess;
  wire                LsuL1Plugin_logic_lsu_ctrl_askRefill;
  wire                LsuL1Plugin_logic_lsu_ctrl_askUpgrade;
  wire                LsuL1Plugin_logic_lsu_ctrl_askFlush;
  wire                LsuL1Plugin_logic_lsu_ctrl_askCbm;
  wire                LsuL1Plugin_logic_lsu_ctrl_doRefill;
  wire                LsuL1Plugin_logic_lsu_ctrl_doUpgrade;
  wire                LsuL1Plugin_logic_lsu_ctrl_doFlush;
  wire                LsuL1Plugin_logic_lsu_ctrl_doWrite;
  wire                LsuL1Plugin_logic_lsu_ctrl_doCbm;
  wire       [0:0]    LsuL1Plugin_logic_lsu_ctrl_wayId;
  wire       [0:0]    LsuL1Plugin_logic_lsu_ctrl_targetWay;
  wire                LsuL1Plugin_logic_lsu_ctrl_doRefillPush;
  wire                when_LsuL1Plugin_l926;
  wire       [2:0]    _zz_22;
  wire                when_LsuL1Plugin_l940;
  wire                when_LsuL1Plugin_l940_1;
  wire       [19:0]   _zz_LsuL1Plugin_logic_waysWrite_tag_address;
  wire                when_LsuL1Plugin_l1028;
  wire                when_LsuL1Plugin_l1035;
  wire                when_LsuL1Plugin_l1039;
  wire                when_LsuL1Plugin_l1039_1;
  wire                when_LsuL1Plugin_l1039_2;
  wire                when_LsuL1Plugin_l1039_3;
  wire                when_LsuL1Plugin_l1039_4;
  wire                when_LsuL1Plugin_l1039_5;
  wire                when_LsuL1Plugin_l1039_6;
  wire                when_LsuL1Plugin_l1039_7;
  wire                when_LsuL1Plugin_l1035_1;
  wire                when_LsuL1Plugin_l1039_8;
  wire                when_LsuL1Plugin_l1039_9;
  wire                when_LsuL1Plugin_l1039_10;
  wire                when_LsuL1Plugin_l1039_11;
  wire                when_LsuL1Plugin_l1039_12;
  wire                when_LsuL1Plugin_l1039_13;
  wire                when_LsuL1Plugin_l1039_14;
  wire                when_LsuL1Plugin_l1039_15;
  reg        [6:0]    LsuL1Plugin_logic_initializer_counter;
  wire                LsuL1Plugin_logic_initializer_done;
  wire                when_LsuL1Plugin_l1233;
  wire       [2:0]    _zz_LsuL1Plugin_logic_shared_write_payload_data_plru_0;
  wire                early0_MulPlugin_logic_formatBus_valid;
  wire       [63:0]   early0_MulPlugin_logic_formatBus_payload;
  reg        [60:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0;
  reg        [60:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_1;
  reg        [60:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_2;
  reg        [60:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_3;
  reg        [60:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_4;
  reg        [60:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_5;
  reg        [60:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_6;
  reg        [43:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0;
  reg        [43:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_1;
  reg        [43:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_2;
  reg        [43:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_3;
  reg        [43:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_4;
  reg        [43:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_5;
  reg        [43:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_6;
  reg        [22:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0;
  reg        [22:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_1;
  reg        [22:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_2;
  reg        [22:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_3;
  reg        [22:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_4;
  reg        [22:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_5;
  reg        [22:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_6;
  reg        [130:0]  _zz_execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0;
  reg        [130:0]  _zz_execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0_1;
  reg                 early0_MulPlugin_logic_writeback_buffer_valid;
  reg        [63:0]   early0_MulPlugin_logic_writeback_buffer_data;
  wire                early0_DivPlugin_logic_formatBus_valid;
  wire       [63:0]   early0_DivPlugin_logic_formatBus_payload;
  reg                 early0_DivPlugin_logic_processing_divRevertResult;
  reg                 early0_DivPlugin_logic_processing_cmdSent;
  wire                io_cmd_fire;
  wire                early0_DivPlugin_logic_processing_request;
  wire       [63:0]   early0_DivPlugin_logic_processing_a;
  wire       [63:0]   early0_DivPlugin_logic_processing_b;
  reg        [63:0]   early0_DivPlugin_logic_processing_a_delay_1;
  reg        [63:0]   early0_DivPlugin_logic_processing_b_delay_1;
  reg                 early0_DivPlugin_logic_processing_relaxer_hadRequest;
  wire                when_DivPlugin_l121;
  reg                 early0_DivPlugin_logic_processing_unscheduleRequest;
  wire                early0_DivPlugin_logic_processing_freeze;
  wire       [63:0]   early0_DivPlugin_logic_processing_selected;
  wire       [63:0]   _zz_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0;
  wire                CsrAccessPlugin_logic_wbWi_valid;
  wire       [63:0]   CsrAccessPlugin_logic_wbWi_payload;
  reg                 CsrAccessPlugin_logic_flushPort_valid;
  reg                 TrapPlugin_logic_fetchL1Invalidate_0_cmd_valid;
  reg                 TrapPlugin_logic_fetchL1Invalidate_0_cmd_ready;
  reg                 TrapPlugin_logic_lsuL1Invalidate_0_cmd_valid;
  wire                TrapPlugin_logic_lsuL1Invalidate_0_cmd_ready;
  reg                 early0_EnvPlugin_logic_trapPort_valid;
  reg                 early0_EnvPlugin_logic_trapPort_payload_exception;
  wire       [38:0]   early0_EnvPlugin_logic_trapPort_payload_tval;
  reg        [3:0]    early0_EnvPlugin_logic_trapPort_payload_code;
  reg        [2:0]    early0_EnvPlugin_logic_trapPort_payload_arg;
  reg                 early0_EnvPlugin_logic_flushPort_valid;
  wire                WhiteboxerPlugin_logic_fetch_fire;
  wire       [38:0]   PrivilegedPlugin_api_lsuTriggerBus_virtual;
  wire       [1:0]    PrivilegedPlugin_api_lsuTriggerBus_size;
  wire                PrivilegedPlugin_api_harts_0_allowInterrupts;
  wire                PrivilegedPlugin_api_harts_0_allowException;
  wire                PrivilegedPlugin_api_harts_0_allowEbreakException;
  wire                PrivilegedPlugin_api_harts_0_fpuEnable;
  wire                LsuL1Plugin_logic_bus_toAxi4_awRaw_valid;
  reg                 LsuL1Plugin_logic_bus_toAxi4_awRaw_ready;
  wire                LsuL1Plugin_logic_bus_toAxi4_awRaw_payload_last;
  wire       [31:0]   LsuL1Plugin_logic_bus_toAxi4_awRaw_payload_fragment_address;
  wire       [63:0]   LsuL1Plugin_logic_bus_toAxi4_awRaw_payload_fragment_data;
  wire                LsuL1Plugin_logic_bus_toAxi4_wRaw_valid;
  wire                LsuL1Plugin_logic_bus_toAxi4_wRaw_ready;
  wire                LsuL1Plugin_logic_bus_toAxi4_wRaw_payload_last;
  wire       [31:0]   LsuL1Plugin_logic_bus_toAxi4_wRaw_payload_fragment_address;
  wire       [63:0]   LsuL1Plugin_logic_bus_toAxi4_wRaw_payload_fragment_data;
  reg                 LsuL1Plugin_logic_bus_write_cmd_fork2_logic_linkEnable_0;
  reg                 LsuL1Plugin_logic_bus_write_cmd_fork2_logic_linkEnable_1;
  wire                when_Stream_l1253;
  wire                when_Stream_l1253_1;
  wire                LsuL1Plugin_logic_bus_toAxi4_awRaw_fire;
  wire                LsuL1Plugin_logic_bus_toAxi4_wRaw_fire;
  reg                 LsuL1Plugin_logic_bus_toAxi4_awRaw_payload_first;
  wire                when_Stream_l581;
  reg                 LsuL1Plugin_logic_bus_toAxi4_awFiltred_valid;
  reg                 LsuL1Plugin_logic_bus_toAxi4_awFiltred_ready;
  wire                LsuL1Plugin_logic_bus_toAxi4_awFiltred_payload_last;
  wire       [31:0]   LsuL1Plugin_logic_bus_toAxi4_awFiltred_payload_fragment_address;
  wire       [63:0]   LsuL1Plugin_logic_bus_toAxi4_awFiltred_payload_fragment_data;
  wire                LsuL1Plugin_logic_bus_toAxi4_aw_valid;
  wire                LsuL1Plugin_logic_bus_toAxi4_aw_ready;
  wire                LsuL1Plugin_logic_bus_toAxi4_aw_payload_last;
  wire       [31:0]   LsuL1Plugin_logic_bus_toAxi4_aw_payload_fragment_address;
  wire       [63:0]   LsuL1Plugin_logic_bus_toAxi4_aw_payload_fragment_data;
  reg                 LsuL1Plugin_logic_bus_toAxi4_awFiltred_rValid;
  reg                 LsuL1Plugin_logic_bus_toAxi4_awFiltred_rData_last;
  reg        [31:0]   LsuL1Plugin_logic_bus_toAxi4_awFiltred_rData_fragment_address;
  reg        [63:0]   LsuL1Plugin_logic_bus_toAxi4_awFiltred_rData_fragment_data;
  wire                when_Stream_l477_1;
  wire                _zz_LsuL1Plugin_logic_bus_toAxi4_wRaw_ready;
  wire                LsuL1Plugin_logic_bus_toAxi4_w_valid;
  wire                LsuL1Plugin_logic_bus_toAxi4_w_ready;
  wire                LsuL1Plugin_logic_bus_toAxi4_w_payload_last;
  wire       [31:0]   LsuL1Plugin_logic_bus_toAxi4_w_payload_fragment_address;
  wire       [63:0]   LsuL1Plugin_logic_bus_toAxi4_w_payload_fragment_data;
  reg        [3:0]    CsrAccessPlugin_bus_decode_trapCode;
  wire                CsrAccessPlugin_bus_decode_fence;
  wire                CsrAccessPlugin_bus_read_valid;
  wire                CsrAccessPlugin_bus_read_moving;
  wire       [11:0]   CsrAccessPlugin_bus_read_address;
  reg                 CsrAccessPlugin_bus_read_halt;
  reg        [63:0]   CsrAccessPlugin_bus_read_toWriteBits;
  wire       [63:0]   CsrAccessPlugin_bus_read_data;
  wire                CsrAccessPlugin_bus_write_valid;
  wire                CsrAccessPlugin_bus_write_moving;
  reg                 CsrAccessPlugin_bus_write_halt;
  reg        [63:0]   CsrAccessPlugin_bus_write_bits;
  wire       [11:0]   CsrAccessPlugin_bus_write_address;
  reg        [3:0]    FetchL1Plugin_logic_trapPort_payload_code;
  reg        [2:0]    FetchL1Plugin_logic_trapPort_payload_arg;
  wire                FetchL1Plugin_logic_events_access;
  wire                FetchL1Plugin_logic_events_miss;
  wire                FetchL1Plugin_logic_events_waiting;
  wire                FetchL1Plugin_logic_banks_0_write_valid;
  wire       [8:0]    FetchL1Plugin_logic_banks_0_write_payload_address;
  wire       [63:0]   FetchL1Plugin_logic_banks_0_write_payload_data;
  wire                FetchL1Plugin_logic_banks_0_read_cmd_valid;
  wire       [8:0]    FetchL1Plugin_logic_banks_0_read_cmd_payload;
  (* keep , syn_keep *) wire       [63:0]   FetchL1Plugin_logic_banks_0_read_rsp /* synthesis syn_keep = 1 */ ;
  wire                FetchL1Plugin_logic_banks_1_write_valid;
  wire       [8:0]    FetchL1Plugin_logic_banks_1_write_payload_address;
  wire       [63:0]   FetchL1Plugin_logic_banks_1_write_payload_data;
  wire                FetchL1Plugin_logic_banks_1_read_cmd_valid;
  wire       [8:0]    FetchL1Plugin_logic_banks_1_read_cmd_payload;
  (* keep , syn_keep *) wire       [63:0]   FetchL1Plugin_logic_banks_1_read_rsp /* synthesis syn_keep = 1 */ ;
  reg        [1:0]    FetchL1Plugin_logic_waysWrite_mask;
  reg        [5:0]    FetchL1Plugin_logic_waysWrite_address;
  reg                 FetchL1Plugin_logic_waysWrite_tag_loaded;
  reg                 FetchL1Plugin_logic_waysWrite_tag_error;
  reg        [19:0]   FetchL1Plugin_logic_waysWrite_tag_address;
  wire                FetchL1Plugin_logic_ways_0_read_cmd_valid;
  wire       [5:0]    FetchL1Plugin_logic_ways_0_read_cmd_payload;
  (* keep , syn_keep *) wire                FetchL1Plugin_logic_ways_0_read_rsp_loaded /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                FetchL1Plugin_logic_ways_0_read_rsp_error /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [19:0]   FetchL1Plugin_logic_ways_0_read_rsp_address /* synthesis syn_keep = 1 */ ;
  wire       [21:0]   _zz_FetchL1Plugin_logic_ways_0_read_rsp_loaded;
  wire                FetchL1Plugin_logic_ways_1_read_cmd_valid;
  wire       [5:0]    FetchL1Plugin_logic_ways_1_read_cmd_payload;
  (* keep , syn_keep *) wire                FetchL1Plugin_logic_ways_1_read_rsp_loaded /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                FetchL1Plugin_logic_ways_1_read_rsp_error /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [19:0]   FetchL1Plugin_logic_ways_1_read_rsp_address /* synthesis syn_keep = 1 */ ;
  wire       [21:0]   _zz_FetchL1Plugin_logic_ways_1_read_rsp_loaded;
  reg                 FetchL1Plugin_logic_plru_write_valid;
  reg        [5:0]    FetchL1Plugin_logic_plru_write_payload_address;
  reg        [0:0]    FetchL1Plugin_logic_plru_write_payload_data_0;
  wire                FetchL1Plugin_logic_plru_read_cmd_valid;
  wire       [5:0]    FetchL1Plugin_logic_plru_read_cmd_payload;
  (* keep , syn_keep *) wire       [0:0]    FetchL1Plugin_logic_plru_read_rsp_0 /* synthesis syn_keep = 1 */ ;
  wire                FetchL1Plugin_logic_invalidate_cmd_valid;
  wire                FetchL1Plugin_logic_invalidate_cmd_ready;
  reg                 FetchL1Plugin_logic_invalidate_canStart;
  reg        [6:0]    FetchL1Plugin_logic_invalidate_counter;
  wire       [6:0]    FetchL1Plugin_logic_invalidate_counterIncr;
  wire                FetchL1Plugin_logic_invalidate_done;
  wire                FetchL1Plugin_logic_invalidate_last;
  reg                 FetchL1Plugin_logic_invalidate_firstEver;
  wire                when_FetchL1Plugin_l204;
  wire                when_FetchL1Plugin_l211;
  wire                when_FetchL1Plugin_l216;
  wire                fetch_logic_ctrls_0_haltRequest_FetchL1Plugin_l217;
  reg                 FetchL1Plugin_logic_refill_start_valid;
  wire       [31:0]   FetchL1Plugin_logic_refill_start_address;
  wire       [0:0]    FetchL1Plugin_logic_refill_start_wayToAllocate;
  wire                FetchL1Plugin_logic_refill_start_isIo;
  reg                 FetchL1Plugin_logic_refill_slots_0_valid;
  reg                 FetchL1Plugin_logic_refill_slots_0_cmdSent;
  (* keep , syn_keep *) reg        [31:0]   FetchL1Plugin_logic_refill_slots_0_address /* synthesis syn_keep = 1 */ ;
  reg                 FetchL1Plugin_logic_refill_slots_0_isIo;
  reg        [0:0]    FetchL1Plugin_logic_refill_slots_0_wayToAllocate;
  reg        [0:0]    FetchL1Plugin_logic_refill_slots_0_priority;
  wire                FetchL1Plugin_logic_refill_slots_0_askCmd;
  reg        [31:0]   FetchL1Plugin_logic_refill_pushCounter;
  wire                FetchL1Plugin_logic_refill_hazard;
  wire                when_FetchL1Plugin_l255;
  wire                when_FetchL1Plugin_l268;
  wire       [0:0]    FetchL1Plugin_logic_refill_onCmd_propoedOh;
  reg                 FetchL1Plugin_logic_refill_onCmd_locked;
  wire                when_FetchL1Plugin_l276;
  reg        [0:0]    FetchL1Plugin_logic_refill_onCmd_lockedOh;
  wire       [0:0]    FetchL1Plugin_logic_refill_onCmd_oh;
  (* keep , syn_keep *) reg        [2:0]    FetchL1Plugin_logic_refill_onRsp_wordIndex /* synthesis syn_keep = 1 */ ;
  wire                FetchL1Plugin_logic_refill_onRsp_holdHarts;
  wire                fetch_logic_ctrls_0_haltRequest_FetchL1Plugin_l297;
  reg                 FetchL1Plugin_logic_refill_onRsp_firstCycle;
  wire                FetchL1Plugin_logic_bus_rsp_fire;
  wire       [0:0]    FetchL1Plugin_logic_refill_onRsp_wayToAllocate;
  wire       [31:0]   FetchL1Plugin_logic_refill_onRsp_address;
  wire                when_FetchL1Plugin_l304;
  wire                when_FetchL1Plugin_l330;
  wire                FetchL1Plugin_logic_cmd_doIt;
  wire                FetchL1Plugin_logic_hits_w_0_indirect_wayTlbHits_0;
  wire                FetchL1Plugin_logic_hits_w_0_indirect_wayTlbHits_1;
  wire                FetchL1Plugin_logic_hits_w_0_indirect_wayTlbHits_2;
  wire                FetchL1Plugin_logic_hits_w_0_indirect_translatedHits;
  wire                FetchL1Plugin_logic_hits_w_0_indirect_bypassHits;
  wire                FetchL1Plugin_logic_hits_w_1_indirect_wayTlbHits_0;
  wire                FetchL1Plugin_logic_hits_w_1_indirect_wayTlbHits_1;
  wire                FetchL1Plugin_logic_hits_w_1_indirect_wayTlbHits_2;
  wire                FetchL1Plugin_logic_hits_w_1_indirect_translatedHits;
  wire                FetchL1Plugin_logic_hits_w_1_indirect_bypassHits;
  wire       [31:0]   FetchL1Plugin_logic_ctrl_pmaPort_cmd_address;
  wire                FetchL1Plugin_logic_ctrl_pmaPort_rsp_fault;
  wire                FetchL1Plugin_logic_ctrl_pmaPort_rsp_io;
  wire       [0:0]    FetchL1Plugin_logic_ctrl_plruLogic_core_io_context_state_0;
  wire       [0:0]    FetchL1Plugin_logic_ctrl_plruLogic_core_io_evict_id;
  wire       [0:0]    FetchL1Plugin_logic_ctrl_plruLogic_core_io_update_id;
  wire       [0:0]    FetchL1Plugin_logic_ctrl_plruLogic_core_io_update_state_0;
  wire                FetchL1Plugin_logic_ctrl_plruLogic_core_evict_sel_0;
  wire                FetchL1Plugin_logic_ctrl_plruLogic_core_evict_logic_0_state;
  wire                FetchL1Plugin_logic_ctrl_plruLogic_buffer_valid;
  wire       [5:0]    FetchL1Plugin_logic_ctrl_plruLogic_buffer_payload_address;
  wire       [0:0]    FetchL1Plugin_logic_ctrl_plruLogic_buffer_payload_data_0;
  reg                 FetchL1Plugin_logic_ctrl_plruLogic_buffer_regNext_valid;
  reg        [5:0]    FetchL1Plugin_logic_ctrl_plruLogic_buffer_regNext_payload_address;
  reg        [0:0]    FetchL1Plugin_logic_ctrl_plruLogic_buffer_regNext_payload_data_0;
  wire                FetchL1Plugin_logic_ctrl_dataAccessFault;
  reg                 FetchL1Plugin_logic_ctrl_trapSent;
  reg                 FetchL1Plugin_logic_ctrl_allowRefill;
  wire                when_FetchL1Plugin_l474;
  wire                when_FetchL1Plugin_l480;
  wire                when_FetchL1Plugin_l487;
  wire                when_FetchL1Plugin_l520;
  wire                when_FetchL1Plugin_l533;
  wire                when_FetchL1Plugin_l537;
  reg                 FetchL1Plugin_logic_ctrl_firstCycle;
  wire                when_FetchL1Plugin_l541;
  reg                 FetchL1Plugin_logic_ctrl_onEvents_waiting;
  wire                when_FetchL1Plugin_l549;
  wire                when_FetchL1Plugin_l558;
  reg        [3:0]    LsuPlugin_logic_trapPort_payload_code;
  reg        [2:0]    LsuPlugin_logic_trapPort_payload_arg;
  reg                 LsuPlugin_logic_flushPort_valid;
  wire       [15:0]   LsuPlugin_logic_flushPort_payload_uopId;
  wire                LsuPlugin_logic_flushPort_payload_self;
  wire                LsuPlugin_logic_frontend_defaultsDecodings_0;
  wire                LsuPlugin_logic_frontend_defaultsDecodings_1;
  wire                LsuPlugin_logic_frontend_defaultsDecodings_2;
  wire                LsuPlugin_logic_frontend_defaultsDecodings_3;
  wire                LsuPlugin_logic_frontend_defaultsDecodings_4;
  wire                LsuPlugin_logic_frontend_defaultsDecodings_5;
  wire                LsuPlugin_logic_commitProbe_valid;
  wire       [38:0]   LsuPlugin_logic_commitProbe_payload_pc;
  wire       [38:0]   LsuPlugin_logic_commitProbe_payload_address;
  wire                LsuPlugin_logic_commitProbe_payload_load;
  wire                LsuPlugin_logic_commitProbe_payload_store;
  wire                LsuPlugin_logic_commitProbe_payload_trap;
  wire                LsuPlugin_logic_commitProbe_payload_io;
  wire                LsuPlugin_logic_commitProbe_payload_prefetchFailed;
  wire                LsuPlugin_logic_commitProbe_payload_miss;
  wire                LsuPlugin_logic_iwb_valid;
  reg        [63:0]   LsuPlugin_logic_iwb_payload;
  reg                 LsuPlugin_logic_cbmCsr_invalIntoClean;
  reg                 PrivilegedPlugin_logic_harts_0_xretAwayFromMachine;
  wire       [0:0]    PrivilegedPlugin_logic_harts_0_commitMask;
  reg                 PrivilegedPlugin_logic_harts_0_int_pending;
  reg        [1:0]    PrivilegedPlugin_logic_harts_0_privilege;
  wire                PrivilegedPlugin_logic_harts_0_withMachinePrivilege;
  wire                PrivilegedPlugin_logic_harts_0_withSupervisorPrivilege;
  wire                PrivilegedPlugin_logic_harts_0_hartRunning;
  wire                PrivilegedPlugin_logic_harts_0_debugMode;
  wire                when_CsrService_l232;
  reg                 PrivilegedPlugin_logic_harts_0_m_status_mie;
  reg                 PrivilegedPlugin_logic_harts_0_m_status_mpie;
  reg        [1:0]    PrivilegedPlugin_logic_harts_0_m_status_mpp;
  reg        [1:0]    PrivilegedPlugin_logic_harts_0_m_status_fs;
  reg                 PrivilegedPlugin_logic_harts_0_m_status_sd;
  reg                 PrivilegedPlugin_logic_harts_0_m_status_tsr;
  reg                 PrivilegedPlugin_logic_harts_0_m_status_tvm;
  reg                 PrivilegedPlugin_logic_harts_0_m_status_tw;
  reg                 PrivilegedPlugin_logic_harts_0_m_status_mprv;
  wire                when_PrivilegedPlugin_l573;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_12;
  wire                when_CsrService_l210;
  reg                 PrivilegedPlugin_logic_harts_0_m_cause_interrupt;
  reg        [3:0]    PrivilegedPlugin_logic_harts_0_m_cause_code;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_13;
  reg                 PrivilegedPlugin_logic_harts_0_m_ip_meip;
  reg                 PrivilegedPlugin_logic_harts_0_m_ip_mtip;
  reg                 PrivilegedPlugin_logic_harts_0_m_ip_msip;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_14;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_15;
  reg                 PrivilegedPlugin_logic_harts_0_m_ie_meie;
  reg                 PrivilegedPlugin_logic_harts_0_m_ie_mtie;
  reg                 PrivilegedPlugin_logic_harts_0_m_ie_msie;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_16;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_17;
  reg                 PrivilegedPlugin_logic_harts_0_m_edeleg_iam;
  reg                 PrivilegedPlugin_logic_harts_0_m_edeleg_bp;
  reg                 PrivilegedPlugin_logic_harts_0_m_edeleg_eu;
  reg                 PrivilegedPlugin_logic_harts_0_m_edeleg_es;
  reg                 PrivilegedPlugin_logic_harts_0_m_edeleg_ipf;
  reg                 PrivilegedPlugin_logic_harts_0_m_edeleg_lpf;
  reg                 PrivilegedPlugin_logic_harts_0_m_edeleg_spf;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_18;
  reg                 PrivilegedPlugin_logic_harts_0_m_ideleg_st;
  reg                 PrivilegedPlugin_logic_harts_0_m_ideleg_se;
  reg                 PrivilegedPlugin_logic_harts_0_m_ideleg_ss;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_19;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_20;
  wire                _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_0_valid;
  wire                _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_1_valid;
  wire                _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_2_valid;
  reg        [3:0]    PrivilegedPlugin_logic_harts_0_m_topi_interrupt;
  wire       [0:0]    PrivilegedPlugin_logic_harts_0_m_topi_priority;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_21;
  reg                 PrivilegedPlugin_logic_harts_0_mcounteren_tm;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_22;
  reg                 PrivilegedPlugin_logic_harts_0_s_cause_interrupt;
  reg        [3:0]    PrivilegedPlugin_logic_harts_0_s_cause_code;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_23;
  reg                 PrivilegedPlugin_logic_harts_0_s_status_sie;
  reg                 PrivilegedPlugin_logic_harts_0_s_status_spie;
  reg        [0:0]    PrivilegedPlugin_logic_harts_0_s_status_spp;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_24;
  reg                 PrivilegedPlugin_logic_harts_0_s_sstc_envcfg_enable;
  wire                PrivilegedPlugin_logic_harts_0_s_sstc_envcfg_allowUpdate;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_25;
  wire                PrivilegedPlugin_logic_harts_0_s_sstc_interrupt;
  reg                 PrivilegedPlugin_logic_harts_0_s_ip_seipSoft;
  reg                 PrivilegedPlugin_logic_harts_0_s_ip_seipInput;
  wire                PrivilegedPlugin_logic_harts_0_s_ip_seipOr;
  reg                 PrivilegedPlugin_logic_harts_0_s_ip_stipSoft;
  wire                PrivilegedPlugin_logic_harts_0_s_ip_stipOr;
  reg                 PrivilegedPlugin_logic_harts_0_s_ip_ssip;
  wire                PrivilegedPlugin_logic_harts_0_s_ip_seipMasked;
  wire                PrivilegedPlugin_logic_harts_0_s_ip_stipMasked;
  wire                PrivilegedPlugin_logic_harts_0_s_ip_ssipMasked;
  reg                 PrivilegedPlugin_logic_harts_0_s_ie_seie;
  reg                 PrivilegedPlugin_logic_harts_0_s_ie_stie;
  reg                 PrivilegedPlugin_logic_harts_0_s_ie_ssie;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_26;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_27;
  wire                when_CsrService_l225;
  wire                _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_0_valid;
  wire                _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_1_valid;
  wire                _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_2_valid;
  reg        [3:0]    PrivilegedPlugin_logic_harts_0_s_topi_interrupt;
  wire       [0:0]    PrivilegedPlugin_logic_harts_0_s_topi_priority;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_28;
  wire                PrivilegedPlugin_logic_harts_0_time_accessable;
  wire       [1:0]    PrivilegedPlugin_logic_defaultTrap_csrPrivilege;
  wire                PrivilegedPlugin_logic_defaultTrap_csrReadOnly;
  wire                when_PrivilegedPlugin_l887;
  wire                GSharePlugin_logic_mem_write_valid;
  wire       [12:0]   GSharePlugin_logic_mem_write_payload_address;
  wire       [1:0]    GSharePlugin_logic_mem_write_payload_data_0;
  wire       [1:0]    GSharePlugin_logic_mem_write_payload_data_1;
  wire                GSharePlugin_logic_mem_writes_0_valid;
  wire       [12:0]   GSharePlugin_logic_mem_writes_0_payload_address;
  wire       [1:0]    GSharePlugin_logic_mem_writes_0_payload_data_0;
  wire       [1:0]    GSharePlugin_logic_mem_writes_0_payload_data_1;
  wire       [12:0]   _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH;
  wire       [12:0]   _zz_GSharePlugin_logic_readRsp_readed_0_0;
  wire       [1:0]    GSharePlugin_logic_readRsp_readed_0_0;
  wire       [1:0]    GSharePlugin_logic_readRsp_readed_0_1;
  wire       [3:0]    _zz_GSharePlugin_logic_readRsp_readed_0_0_1;
  wire                when_GSharePlugin_l100;
  reg        [1:0]    BtbPlugin_logic_ras_ptr_push;
  reg        [1:0]    BtbPlugin_logic_ras_ptr_pop;
  reg                 BtbPlugin_logic_ras_ptr_pushIt;
  reg                 BtbPlugin_logic_ras_ptr_popIt;
  wire                BtbPlugin_logic_ras_readIt;
  reg        [37:0]   BtbPlugin_logic_ras_read;
  wire                BtbPlugin_logic_ras_write_valid;
  wire       [1:0]    BtbPlugin_logic_ras_write_payload_address;
  reg        [37:0]   BtbPlugin_logic_ras_write_payload_data;
  reg                 BtbPlugin_logic_memWrite_valid;
  reg        [8:0]    BtbPlugin_logic_memWrite_payload_address;
  reg        [15:0]   BtbPlugin_logic_memWrite_payload_data_0_hash;
  reg        [0:0]    BtbPlugin_logic_memWrite_payload_data_0_sliceLow;
  wire       [37:0]   BtbPlugin_logic_memWrite_payload_data_0_pcTarget;
  reg                 BtbPlugin_logic_memWrite_payload_data_0_isBranch;
  reg                 BtbPlugin_logic_memWrite_payload_data_0_isPush;
  reg                 BtbPlugin_logic_memWrite_payload_data_0_isPop;
  reg        [0:0]    BtbPlugin_logic_memWrite_payload_mask;
  wire                BtbPlugin_logic_memRead_cmd_valid;
  wire       [8:0]    BtbPlugin_logic_memRead_cmd_payload;
  wire       [15:0]   BtbPlugin_logic_memRead_rsp_0_hash;
  wire       [0:0]    BtbPlugin_logic_memRead_rsp_0_sliceLow;
  wire       [37:0]   BtbPlugin_logic_memRead_rsp_0_pcTarget;
  wire                BtbPlugin_logic_memRead_rsp_0_isBranch;
  wire                BtbPlugin_logic_memRead_rsp_0_isPush;
  wire                BtbPlugin_logic_memRead_rsp_0_isPop;
  wire                BtbPlugin_logic_memDp_wp_valid;
  wire       [8:0]    BtbPlugin_logic_memDp_wp_payload_address;
  wire       [15:0]   BtbPlugin_logic_memDp_wp_payload_data_0_hash;
  wire       [0:0]    BtbPlugin_logic_memDp_wp_payload_data_0_sliceLow;
  wire       [37:0]   BtbPlugin_logic_memDp_wp_payload_data_0_pcTarget;
  wire                BtbPlugin_logic_memDp_wp_payload_data_0_isBranch;
  wire                BtbPlugin_logic_memDp_wp_payload_data_0_isPush;
  wire                BtbPlugin_logic_memDp_wp_payload_data_0_isPop;
  wire       [0:0]    BtbPlugin_logic_memDp_wp_payload_mask;
  wire                BtbPlugin_logic_memDp_rp_cmd_valid;
  wire       [8:0]    BtbPlugin_logic_memDp_rp_cmd_payload;
  wire       [15:0]   BtbPlugin_logic_memDp_rp_rsp_0_hash;
  wire       [0:0]    BtbPlugin_logic_memDp_rp_rsp_0_sliceLow;
  wire       [37:0]   BtbPlugin_logic_memDp_rp_rsp_0_pcTarget;
  wire                BtbPlugin_logic_memDp_rp_rsp_0_isBranch;
  wire                BtbPlugin_logic_memDp_rp_rsp_0_isPush;
  wire                BtbPlugin_logic_memDp_rp_rsp_0_isPop;
  wire       [57:0]   _zz_BtbPlugin_logic_memDp_rp_rsp_0_hash;
  wire       [9:0]    WhiteboxerPlugin_logic_fetch_fetchId;
  wire                WhiteboxerPlugin_logic_decodes_0_fire;
  reg                 decode_ctrls_0_up_LANE_SEL_0_regNext;
  wire                when_CtrlLaneApi_l50;
  wire                WhiteboxerPlugin_logic_decodes_0_spawn;
  wire       [63:0]   WhiteboxerPlugin_logic_decodes_0_pc;
  wire       [9:0]    WhiteboxerPlugin_logic_decodes_0_fetchId;
  wire       [9:0]    WhiteboxerPlugin_logic_decodes_0_decodeId;
  wire       [15:0]   early0_BranchPlugin_logic_flushPort_payload_uopId;
  wire                early0_BranchPlugin_logic_flushPort_payload_self;
  wire       [15:0]   CsrAccessPlugin_logic_flushPort_payload_uopId;
  wire                CsrAccessPlugin_logic_flushPort_payload_self;
  reg                 CsrAccessPlugin_logic_trapPort_valid;
  reg                 CsrAccessPlugin_logic_trapPort_payload_exception;
  wire       [38:0]   CsrAccessPlugin_logic_trapPort_payload_tval;
  reg        [3:0]    CsrAccessPlugin_logic_trapPort_payload_code;
  wire       [2:0]    CsrAccessPlugin_logic_trapPort_payload_arg;
  wire       [15:0]   early0_EnvPlugin_logic_flushPort_payload_uopId;
  wire                early0_EnvPlugin_logic_flushPort_payload_self;
  wire       [3:0]    MmuPlugin_logic_satpModeWrite;
  wire       [31:0]   FetchL1Plugin_pmaBuilder_addressBits;
  wire                _zz_FetchL1Plugin_logic_ctrl_pmaPort_rsp_io;
  wire                FetchL1Plugin_pmaBuilder_onTransfers_0_addressHit;
  wire                FetchL1Plugin_pmaBuilder_onTransfers_0_argsHit;
  wire                FetchL1Plugin_pmaBuilder_onTransfers_0_hit;
  reg                 DecoderPlugin_logic_forgetPort_valid;
  reg        [38:0]   DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice;
  wire       [0:0]    PerformanceCounterPlugin_logic_commitMask;
  reg                 PerformanceCounterPlugin_logic_ignoreNextCommit;
  wire                when_PerformanceCounterPlugin_l45;
  wire       [0:0]    PerformanceCounterPlugin_logic_commitCount;
  wire                PerformanceCounterPlugin_logic_eventCycles;
  wire                PerformanceCounterPlugin_logic_eventInstructions_0;
  reg        [7:0]    PerformanceCounterPlugin_logic_counters_cycle_value;
  wire                PerformanceCounterPlugin_logic_counters_cycle_needFlush;
  reg                 PerformanceCounterPlugin_logic_counters_cycle_mcounteren;
  reg                 PerformanceCounterPlugin_logic_counters_cycle_scounteren;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_29;
  reg                 PerformanceCounterPlugin_logic_counters_cycle_mcountinhibit;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_30;
  reg        [7:0]    PerformanceCounterPlugin_logic_counters_instret_value;
  wire                PerformanceCounterPlugin_logic_counters_instret_needFlush;
  reg                 PerformanceCounterPlugin_logic_counters_instret_mcounteren;
  reg                 PerformanceCounterPlugin_logic_counters_instret_scounteren;
  reg                 PerformanceCounterPlugin_logic_counters_instret_mcountinhibit;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_counters_instret_value;
  wire                LsuPlugin_logic_cbmCsr_menvcfg_privLower;
  reg        [1:0]    LsuPlugin_logic_cbmCsr_menvcfg_cbie;
  reg        [0:0]    LsuPlugin_logic_cbmCsr_menvcfg_cbcfe;
  wire                when_LsuPlugin_l226;
  wire                LsuPlugin_logic_cbmCsr_senvcfg_privLower;
  reg        [1:0]    LsuPlugin_logic_cbmCsr_senvcfg_cbie;
  reg        [0:0]    LsuPlugin_logic_cbmCsr_senvcfg_cbcfe;
  wire                when_LsuPlugin_l226_1;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_31;
  wire                execute_lane0_ctrls_0_upIsCancel;
  wire                execute_lane0_ctrls_0_downIsCancel;
  wire                LsuPlugin_logic_bus_cmd_valid;
  wire                LsuPlugin_logic_bus_cmd_ready;
  wire                LsuPlugin_logic_bus_cmd_payload_write;
  wire       [31:0]   LsuPlugin_logic_bus_cmd_payload_address;
  wire       [63:0]   LsuPlugin_logic_bus_cmd_payload_data;
  wire       [1:0]    LsuPlugin_logic_bus_cmd_payload_size;
  wire       [7:0]    LsuPlugin_logic_bus_cmd_payload_mask;
  wire                LsuPlugin_logic_bus_cmd_payload_io;
  wire                LsuPlugin_logic_bus_cmd_payload_fromHart;
  wire       [15:0]   LsuPlugin_logic_bus_cmd_payload_uopId;
  reg                 LsuPlugin_logic_bus_rsp_valid;
  reg                 LsuPlugin_logic_bus_rsp_payload_error;
  wire       [63:0]   LsuPlugin_logic_bus_rsp_payload_data;
  wire                LsuPlugin_logic_flusher_wantExit;
  reg                 LsuPlugin_logic_flusher_wantStart;
  wire                LsuPlugin_logic_flusher_wantKill;
  reg        [6:0]    LsuPlugin_logic_flusher_cmdCounter;
  wire                LsuPlugin_logic_flusher_inflight;
  reg        [0:0]    LsuPlugin_logic_flusher_waiter;
  wire       [4:0]    LsuPlugin_logic_onAddress0_ls_prefetchOp;
  wire                LsuPlugin_logic_onAddress0_ls_port_valid;
  wire                LsuPlugin_logic_onAddress0_ls_port_ready;
  wire       [2:0]    LsuPlugin_logic_onAddress0_ls_port_payload_op;
  wire       [38:0]   LsuPlugin_logic_onAddress0_ls_port_payload_address;
  wire       [1:0]    LsuPlugin_logic_onAddress0_ls_port_payload_size;
  wire                LsuPlugin_logic_onAddress0_ls_port_payload_load;
  wire                LsuPlugin_logic_onAddress0_ls_port_payload_store;
  wire                LsuPlugin_logic_onAddress0_ls_port_payload_atomic;
  wire                LsuPlugin_logic_onAddress0_ls_port_payload_clean;
  wire                LsuPlugin_logic_onAddress0_ls_port_payload_invalidate;
  wire       [11:0]   LsuPlugin_logic_onAddress0_ls_port_payload_storeId;
  reg        [11:0]   LsuPlugin_logic_onAddress0_ls_storeId;
  wire                LsuPlugin_logic_onAddress0_ls_port_fire;
  reg        [0:0]    LsuPlugin_logic_onAddress0_access_waiter_refill;
  reg                 LsuPlugin_logic_onAddress0_access_waiter_valid;
  wire                when_LsuPlugin_l264;
  wire                LsuPlugin_logic_onAddress0_access_sbWaiter;
  wire                LsuPlugin_logic_onAddress0_access_port_valid;
  wire                LsuPlugin_logic_onAddress0_access_port_ready;
  wire       [2:0]    LsuPlugin_logic_onAddress0_access_port_payload_op;
  wire       [38:0]   LsuPlugin_logic_onAddress0_access_port_payload_address;
  wire       [1:0]    LsuPlugin_logic_onAddress0_access_port_payload_size;
  wire                LsuPlugin_logic_onAddress0_access_port_payload_load;
  wire                LsuPlugin_logic_onAddress0_access_port_payload_store;
  wire                LsuPlugin_logic_onAddress0_access_port_payload_atomic;
  wire                LsuPlugin_logic_onAddress0_access_port_payload_clean;
  wire                LsuPlugin_logic_onAddress0_access_port_payload_invalidate;
  wire       [11:0]   LsuPlugin_logic_onAddress0_access_port_payload_storeId;
  wire                _zz_MmuPlugin_logic_accessBus_cmd_ready;
  wire                MmuPlugin_logic_accessBus_cmd_haltWhen_valid;
  wire                MmuPlugin_logic_accessBus_cmd_haltWhen_ready;
  wire       [31:0]   MmuPlugin_logic_accessBus_cmd_haltWhen_payload_address;
  wire       [1:0]    MmuPlugin_logic_accessBus_cmd_haltWhen_payload_size;
  wire                LsuPlugin_logic_onAddress0_flush_port_valid;
  wire                LsuPlugin_logic_onAddress0_flush_port_ready;
  wire       [2:0]    LsuPlugin_logic_onAddress0_flush_port_payload_op;
  wire       [38:0]   LsuPlugin_logic_onAddress0_flush_port_payload_address;
  wire       [1:0]    LsuPlugin_logic_onAddress0_flush_port_payload_size;
  wire                LsuPlugin_logic_onAddress0_flush_port_payload_load;
  wire                LsuPlugin_logic_onAddress0_flush_port_payload_store;
  wire                LsuPlugin_logic_onAddress0_flush_port_payload_atomic;
  wire                LsuPlugin_logic_onAddress0_flush_port_payload_clean;
  wire                LsuPlugin_logic_onAddress0_flush_port_payload_invalidate;
  wire       [11:0]   LsuPlugin_logic_onAddress0_flush_port_payload_storeId;
  wire                LsuPlugin_logic_onAddress0_flush_port_fire;
  reg        [7:0]    _zz_execute_ctrl2_down_LsuL1_MASK_lane0;
  wire                when_LsuPlugin_l529;
  wire                when_LsuPlugin_l557;
  wire                when_LsuPlugin_l557_1;
  wire                when_LsuPlugin_l565;
  wire       [31:0]   LsuPlugin_logic_onPma_cached_cmd_address;
  wire       [0:0]    LsuPlugin_logic_onPma_cached_cmd_op;
  wire                LsuPlugin_logic_onPma_cached_rsp_fault;
  wire                LsuPlugin_logic_onPma_cached_rsp_io;
  wire       [31:0]   LsuPlugin_logic_onPma_io_cmd_address;
  wire       [1:0]    LsuPlugin_logic_onPma_io_cmd_size;
  wire       [0:0]    LsuPlugin_logic_onPma_io_cmd_op;
  wire                LsuPlugin_logic_onPma_io_rsp_fault;
  wire                LsuPlugin_logic_onPma_io_rsp_io;
  wire                when_LsuPlugin_l580;
  wire                LsuPlugin_logic_onPma_addressExtension;
  wire       [24:0]   _zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0;
  reg                 LsuPlugin_logic_onCtrl_lsuTrap;
  reg        [63:0]   LsuPlugin_logic_onCtrl_writeData;
  wire                LsuPlugin_logic_onCtrl_scMiss;
  reg                 LsuPlugin_logic_onCtrl_io_tooEarly;
  reg                 LsuPlugin_logic_onCtrl_io_allowIt;
  wire                when_LsuPlugin_l608;
  wire                LsuPlugin_logic_onCtrl_io_doIt;
  reg                 LsuPlugin_logic_onCtrl_io_doItReg;
  reg                 LsuPlugin_logic_onCtrl_io_cmdSent;
  wire                LsuPlugin_logic_bus_cmd_fire;
  wire                when_LsuPlugin_l612;
  wire                LsuPlugin_logic_bus_rsp_toStream_valid;
  wire                LsuPlugin_logic_bus_rsp_toStream_ready;
  wire                LsuPlugin_logic_bus_rsp_toStream_payload_error;
  wire       [63:0]   LsuPlugin_logic_bus_rsp_toStream_payload_data;
  wire                LsuPlugin_logic_onCtrl_io_rsp_valid;
  wire                LsuPlugin_logic_onCtrl_io_rsp_ready;
  wire                LsuPlugin_logic_onCtrl_io_rsp_payload_error;
  wire       [63:0]   LsuPlugin_logic_onCtrl_io_rsp_payload_data;
  reg                 LsuPlugin_logic_bus_rsp_toStream_rValid;
  wire                LsuPlugin_logic_onCtrl_io_rsp_fire;
  reg                 LsuPlugin_logic_bus_rsp_toStream_rData_error;
  reg        [63:0]   LsuPlugin_logic_bus_rsp_toStream_rData_data;
  wire                LsuPlugin_logic_onCtrl_io_freezeIt;
  wire       [63:0]   LsuPlugin_logic_onCtrl_loadData_input;
  wire       [7:0]    LsuPlugin_logic_onCtrl_loadData_splitted_0;
  wire       [7:0]    LsuPlugin_logic_onCtrl_loadData_splitted_1;
  wire       [7:0]    LsuPlugin_logic_onCtrl_loadData_splitted_2;
  wire       [7:0]    LsuPlugin_logic_onCtrl_loadData_splitted_3;
  wire       [7:0]    LsuPlugin_logic_onCtrl_loadData_splitted_4;
  wire       [7:0]    LsuPlugin_logic_onCtrl_loadData_splitted_5;
  wire       [7:0]    LsuPlugin_logic_onCtrl_loadData_splitted_6;
  wire       [7:0]    LsuPlugin_logic_onCtrl_loadData_splitted_7;
  reg        [63:0]   LsuPlugin_logic_onCtrl_loadData_shifted;
  wire       [63:0]   LsuPlugin_logic_onCtrl_storeData_mapping_0_1;
  wire       [63:0]   LsuPlugin_logic_onCtrl_storeData_mapping_1_1;
  wire       [63:0]   LsuPlugin_logic_onCtrl_storeData_mapping_2_1;
  wire       [63:0]   LsuPlugin_logic_onCtrl_storeData_mapping_3_1;
  reg        [63:0]   _zz_execute_ctrl4_down_LsuL1_WRITE_DATA_lane0;
  reg        [63:0]   LsuPlugin_logic_onCtrl_rva_srcBuffer;
  wire       [2:0]    _zz_LsuPlugin_logic_onCtrl_rva_alu_compare;
  wire                _zz_LsuPlugin_logic_onCtrl_rva_alu_selectRf;
  wire                when_Rvi_l230;
  wire                LsuPlugin_logic_onCtrl_rva_alu_compare;
  wire                LsuPlugin_logic_onCtrl_rva_alu_unsigned;
  wire       [63:0]   LsuPlugin_logic_onCtrl_rva_alu_addSub;
  reg                 LsuPlugin_logic_onCtrl_rva_alu_less;
  wire                LsuPlugin_logic_onCtrl_rva_alu_selectRf;
  wire       [2:0]    switch_Misc_l245;
  reg        [63:0]   LsuPlugin_logic_onCtrl_rva_alu_raw;
  reg        [63:0]   LsuPlugin_logic_onCtrl_rva_alu_result;
  reg        [63:0]   LsuPlugin_logic_onCtrl_rva_aluBuffer;
  wire                LsuPlugin_logic_onCtrl_rva_delay_0;
  wire                LsuPlugin_logic_onCtrl_rva_delay_1;
  reg                 _zz_LsuPlugin_logic_onCtrl_rva_delay_0;
  reg                 _zz_LsuPlugin_logic_onCtrl_rva_delay_1;
  wire                LsuPlugin_logic_onCtrl_rva_freezeIt;
  reg                 LsuPlugin_logic_onCtrl_rva_lrsc_capture;
  reg                 LsuPlugin_logic_onCtrl_rva_lrsc_reserved;
  reg        [31:0]   LsuPlugin_logic_onCtrl_rva_lrsc_address;
  wire                when_LsuPlugin_l697;
  reg        [5:0]    LsuPlugin_logic_onCtrl_rva_lrsc_age;
  wire                when_LsuPlugin_l709;
  wire                when_LsuPlugin_l716;
  wire                when_LsuPlugin_l720;
  wire                LsuPlugin_logic_onCtrl_traps_accessFault;
  wire                LsuPlugin_logic_onCtrl_traps_l1Failed;
  wire                LsuPlugin_logic_onCtrl_traps_pmaFault;
  wire                when_LsuPlugin_l820;
  wire                when_LsuPlugin_l847;
  wire                LsuPlugin_logic_onCtrl_fenceTrap_enable;
  reg                 LsuPlugin_logic_onCtrl_fenceTrap_doIt;
  reg                 LsuPlugin_logic_onCtrl_fenceTrap_doItReg;
  wire                when_LsuPlugin_l855;
  wire                when_LsuPlugin_l857;
  wire                when_LsuPlugin_l897;
  reg                 LsuPlugin_logic_onCtrl_cmbTrap_cmbTrigger;
  reg        [0:0]    LsuPlugin_logic_onCtrl_cmbTrap_pendingWritebacks;
  wire                LsuPlugin_logic_onCtrl_cmbTrap_pending;
  wire                LsuPlugin_logic_onCtrl_cmbTrap_valid;
  wire                when_LsuPlugin_l908;
  wire                LsuPlugin_logic_onCtrl_mmuNeeded;
  wire                when_LsuPlugin_l949;
  wire                when_LsuPlugin_l986;
  wire                when_LsuPlugin_l268;
  reg        [0:0]    LsuPlugin_logic_onCtrl_hartRegulation_refill;
  reg                 LsuPlugin_logic_onCtrl_hartRegulation_valid;
  wire                when_LsuPlugin_l264_1;
  wire                when_LsuPlugin_l993;
  wire                when_LsuPlugin_l268_1;
  wire                LsuPlugin_logic_onCtrl_commitProbeReq;
  reg                 LsuPlugin_logic_onCtrl_commitProbeToken;
  wire                when_LsuPlugin_l1018;
  wire                LsuPlugin_logic_onWb_storeFire;
  wire                LsuPlugin_logic_onWb_storeBroadcast;
  wire                execute_lane0_ctrls_1_upIsCancel;
  wire                execute_lane0_ctrls_1_downIsCancel;
  reg        [63:0]   _zz_execute_ctrl1_down_early0_SrcPlugin_SRC1_lane0;
  reg        [63:0]   _zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0;
  reg        [63:0]   early0_SrcPlugin_logic_addsub_combined_rs2Patched;
  wire                lane0_IntFormatPlugin_logic_stages_0_wb_valid;
  reg        [63:0]   lane0_IntFormatPlugin_logic_stages_0_wb_payload;
  wire       [1:0]    lane0_IntFormatPlugin_logic_stages_0_hits;
  wire       [63:0]   lane0_IntFormatPlugin_logic_stages_0_raw;
  wire                lane0_IntFormatPlugin_logic_stages_0_segments_0_sign_sels_0;
  reg                 _zz_lane0_IntFormatPlugin_logic_stages_0_segments_0_sign_value;
  wire                lane0_IntFormatPlugin_logic_stages_0_segments_0_sign_value;
  wire                lane0_IntFormatPlugin_logic_stages_0_segments_0_doIt;
  wire                lane0_IntFormatPlugin_logic_stages_1_wb_valid;
  reg        [63:0]   lane0_IntFormatPlugin_logic_stages_1_wb_payload;
  wire       [1:0]    lane0_IntFormatPlugin_logic_stages_1_hits;
  wire       [63:0]   lane0_IntFormatPlugin_logic_stages_1_raw;
  wire                lane0_IntFormatPlugin_logic_stages_1_segments_0_sign_sels_0;
  reg                 _zz_lane0_IntFormatPlugin_logic_stages_1_segments_0_sign_value;
  wire                lane0_IntFormatPlugin_logic_stages_1_segments_0_sign_value;
  wire                lane0_IntFormatPlugin_logic_stages_1_segments_0_doIt;
  wire                lane0_IntFormatPlugin_logic_stages_1_segments_1_sign_sels_0;
  wire                lane0_IntFormatPlugin_logic_stages_1_segments_1_sign_sels_1;
  reg                 _zz_lane0_IntFormatPlugin_logic_stages_1_segments_1_sign_value;
  wire                lane0_IntFormatPlugin_logic_stages_1_segments_1_sign_value;
  wire                lane0_IntFormatPlugin_logic_stages_1_segments_1_doIt;
  wire                lane0_IntFormatPlugin_logic_stages_1_segments_2_sign_sels_0;
  wire                lane0_IntFormatPlugin_logic_stages_1_segments_2_sign_sels_1;
  wire                lane0_IntFormatPlugin_logic_stages_1_segments_2_sign_sels_2;
  reg                 _zz_lane0_IntFormatPlugin_logic_stages_1_segments_2_sign_value;
  wire                lane0_IntFormatPlugin_logic_stages_1_segments_2_sign_value;
  wire                lane0_IntFormatPlugin_logic_stages_1_segments_2_doIt;
  wire                lane0_IntFormatPlugin_logic_stages_2_wb_valid;
  reg        [63:0]   lane0_IntFormatPlugin_logic_stages_2_wb_payload;
  wire       [1:0]    lane0_IntFormatPlugin_logic_stages_2_hits;
  wire       [63:0]   lane0_IntFormatPlugin_logic_stages_2_raw;
  wire                lane0_IntFormatPlugin_logic_stages_2_segments_0_sign_sels_0;
  reg                 _zz_lane0_IntFormatPlugin_logic_stages_2_segments_0_sign_value;
  wire                lane0_IntFormatPlugin_logic_stages_2_segments_0_sign_value;
  wire                lane0_IntFormatPlugin_logic_stages_2_segments_0_doIt;
  reg        [38:0]   early0_BranchPlugin_pcCalc_target_a;
  reg        [63:0]   early0_BranchPlugin_pcCalc_target_b;
  wire       [1:0]    early0_BranchPlugin_pcCalc_slices;
  wire       [1:0]    AlignerPlugin_logic_maskGen_frontMasks_0;
  wire       [1:0]    AlignerPlugin_logic_maskGen_frontMasks_1;
  wire       [1:0]    AlignerPlugin_logic_maskGen_backMasks_0;
  wire       [1:0]    AlignerPlugin_logic_maskGen_backMasks_1;
  wire       [15:0]   AlignerPlugin_logic_slices_data_0;
  wire       [15:0]   AlignerPlugin_logic_slices_data_1;
  wire       [15:0]   AlignerPlugin_logic_slices_data_2;
  wire       [15:0]   AlignerPlugin_logic_slices_data_3;
  wire       [3:0]    AlignerPlugin_logic_slices_mask;
  wire       [3:0]    AlignerPlugin_logic_slices_last;
  wire       [31:0]   AlignerPlugin_logic_slicesInstructions_0;
  wire       [31:0]   AlignerPlugin_logic_slicesInstructions_1;
  wire       [31:0]   AlignerPlugin_logic_slicesInstructions_2;
  wire       [31:0]   AlignerPlugin_logic_slicesInstructions_3;
  reg        [3:0]    AlignerPlugin_logic_scanners_0_usageMask;
  wire                AlignerPlugin_logic_scanners_0_checker_0_required;
  wire                AlignerPlugin_logic_scanners_0_checker_0_last;
  wire                AlignerPlugin_logic_scanners_0_checker_0_redo;
  wire                AlignerPlugin_logic_scanners_0_checker_0_present;
  wire                AlignerPlugin_logic_scanners_0_checker_0_valid;
  wire                AlignerPlugin_logic_scanners_0_checker_1_required;
  wire                AlignerPlugin_logic_scanners_0_checker_1_last;
  wire                AlignerPlugin_logic_scanners_0_checker_1_redo;
  wire                AlignerPlugin_logic_scanners_0_checker_1_present;
  wire                AlignerPlugin_logic_scanners_0_checker_1_valid;
  wire                AlignerPlugin_logic_scanners_0_redo;
  wire                AlignerPlugin_logic_scanners_0_valid;
  reg        [3:0]    AlignerPlugin_logic_scanners_1_usageMask;
  wire                AlignerPlugin_logic_scanners_1_checker_0_required;
  wire                AlignerPlugin_logic_scanners_1_checker_0_last;
  wire                AlignerPlugin_logic_scanners_1_checker_0_redo;
  wire                AlignerPlugin_logic_scanners_1_checker_0_present;
  wire                AlignerPlugin_logic_scanners_1_checker_0_valid;
  wire                AlignerPlugin_logic_scanners_1_checker_1_required;
  wire                AlignerPlugin_logic_scanners_1_checker_1_last;
  wire                AlignerPlugin_logic_scanners_1_checker_1_redo;
  wire                AlignerPlugin_logic_scanners_1_checker_1_present;
  wire                AlignerPlugin_logic_scanners_1_checker_1_valid;
  wire                AlignerPlugin_logic_scanners_1_redo;
  wire                AlignerPlugin_logic_scanners_1_valid;
  reg        [3:0]    AlignerPlugin_logic_scanners_2_usageMask;
  wire                AlignerPlugin_logic_scanners_2_checker_0_required;
  wire                AlignerPlugin_logic_scanners_2_checker_0_last;
  wire                AlignerPlugin_logic_scanners_2_checker_0_redo;
  wire                AlignerPlugin_logic_scanners_2_checker_0_present;
  wire                AlignerPlugin_logic_scanners_2_checker_0_valid;
  wire                AlignerPlugin_logic_scanners_2_checker_1_required;
  wire                AlignerPlugin_logic_scanners_2_checker_1_last;
  wire                AlignerPlugin_logic_scanners_2_checker_1_redo;
  wire                AlignerPlugin_logic_scanners_2_checker_1_present;
  wire                AlignerPlugin_logic_scanners_2_checker_1_valid;
  wire                AlignerPlugin_logic_scanners_2_redo;
  wire                AlignerPlugin_logic_scanners_2_valid;
  reg        [3:0]    AlignerPlugin_logic_scanners_3_usageMask;
  wire                AlignerPlugin_logic_scanners_3_checker_0_required;
  wire                AlignerPlugin_logic_scanners_3_checker_0_last;
  wire                AlignerPlugin_logic_scanners_3_checker_0_redo;
  wire                AlignerPlugin_logic_scanners_3_checker_0_present;
  wire                AlignerPlugin_logic_scanners_3_checker_0_valid;
  wire                AlignerPlugin_logic_scanners_3_checker_1_required;
  wire                AlignerPlugin_logic_scanners_3_checker_1_last;
  wire                AlignerPlugin_logic_scanners_3_checker_1_redo;
  wire                AlignerPlugin_logic_scanners_3_checker_1_present;
  wire                AlignerPlugin_logic_scanners_3_checker_1_valid;
  wire                AlignerPlugin_logic_scanners_3_redo;
  wire                AlignerPlugin_logic_scanners_3_valid;
  wire       [3:0]    AlignerPlugin_logic_usedMask_0;
  wire       [3:0]    AlignerPlugin_logic_usedMask_1;
  wire                AlignerPlugin_logic_extractors_0_first;
  wire       [3:0]    AlignerPlugin_logic_extractors_0_usableMask;
  wire       [3:0]    _zz_AlignerPlugin_logic_extractors_0_usableMask_bools_0;
  wire                AlignerPlugin_logic_extractors_0_usableMask_bools_0;
  wire                AlignerPlugin_logic_extractors_0_usableMask_bools_1;
  wire                AlignerPlugin_logic_extractors_0_usableMask_bools_2;
  wire                AlignerPlugin_logic_extractors_0_usableMask_bools_3;
  reg        [3:0]    _zz_AlignerPlugin_logic_extractors_0_slicesOh;
  wire                AlignerPlugin_logic_extractors_0_usableMask_range_0_to_1;
  wire                AlignerPlugin_logic_extractors_0_usableMask_range_0_to_2;
  wire       [3:0]    AlignerPlugin_logic_extractors_0_slicesOh;
  wire                _zz_AlignerPlugin_logic_extractors_0_redo;
  wire                _zz_AlignerPlugin_logic_extractors_0_redo_1;
  wire                _zz_AlignerPlugin_logic_extractors_0_redo_2;
  wire                _zz_AlignerPlugin_logic_extractors_0_redo_3;
  reg                 AlignerPlugin_logic_extractors_0_redo;
  wire       [1:0]    AlignerPlugin_logic_extractors_0_localMask;
  wire       [3:0]    AlignerPlugin_logic_extractors_0_usageMask;
  reg                 AlignerPlugin_logic_extractors_0_valid;
  reg        [38:0]   AlignerPlugin_logic_extractors_0_ctx_pc;
  wire       [31:0]   AlignerPlugin_logic_extractors_0_ctx_instruction;
  wire       [9:0]    AlignerPlugin_logic_extractors_0_ctx_hm_Fetch_ID;
  wire       [1:0]    AlignerPlugin_logic_extractors_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    AlignerPlugin_logic_extractors_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_1;
  wire       [11:0]   AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_BRANCH_HISTORY;
  wire       [1:0]    AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_SLICES_BRANCH;
  wire       [1:0]    AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_SLICES_TAKEN;
  wire       [38:0]   AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_JUMP_PC;
  wire                AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_JUMPED;
  wire       [0:0]    AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_JUMP_SLICE;
  wire                AlignerPlugin_logic_extractors_0_ctx_trap;
  wire                when_AlignerPlugin_l160;
  reg        [9:0]    AlignerPlugin_logic_feeder_harts_0_dopId;
  wire                when_AlignerPlugin_l171;
  wire                AlignerPlugin_logic_feeder_lanes_0_valid;
  wire                AlignerPlugin_logic_feeder_lanes_0_isRvc;
  reg        [31:0]   AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst;
  reg                 AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_illegal;
  wire       [4:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst;
  wire       [4:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_1;
  wire       [11:0]   _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_2;
  wire       [11:0]   _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_3;
  wire                _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_4;
  reg        [11:0]   _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_5;
  wire                _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_6;
  reg        [14:0]   _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_7;
  wire                _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_8;
  reg        [2:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_9;
  wire                _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10;
  reg        [9:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_11;
  wire       [20:0]   _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_12;
  wire                _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_13;
  reg        [4:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_14;
  wire       [12:0]   _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_15;
  wire       [4:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_16;
  wire       [4:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_17;
  wire       [4:0]    switch_Rvc_l55;
  wire                when_Rvc_l59;
  wire                when_Rvc_l73;
  wire                when_Rvc_l80;
  wire       [31:0]   _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_18;
  wire                when_Rvc_l101;
  wire                when_Rvc_l106;
  wire                when_Rvc_l114;
  wire       [1:0]    _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0;
  wire       [1:0]    _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_1;
  wire                _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_2;
  reg        [1:0]    _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_3;
  wire       [1:0]    _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_4;
  wire                _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_5;
  wire       [0:0]    AlignerPlugin_logic_feeder_lanes_0_onBtb_pcLastSlice;
  wire                AlignerPlugin_logic_feeder_lanes_0_onBtb_didPrediction;
  reg        [31:0]   AlignerPlugin_logic_buffer_data;
  reg        [1:0]    AlignerPlugin_logic_buffer_mask;
  reg        [1:0]    AlignerPlugin_logic_buffer_last;
  reg        [38:0]   AlignerPlugin_logic_buffer_pc;
  reg                 AlignerPlugin_logic_buffer_trap;
  reg        [9:0]    AlignerPlugin_logic_buffer_hm_Fetch_ID;
  reg        [1:0]    AlignerPlugin_logic_buffer_hm_GSharePlugin_GSHARE_COUNTER_0;
  reg        [1:0]    AlignerPlugin_logic_buffer_hm_GSharePlugin_GSHARE_COUNTER_1;
  reg        [11:0]   AlignerPlugin_logic_buffer_hm_Prediction_BRANCH_HISTORY;
  reg        [1:0]    AlignerPlugin_logic_buffer_hm_Prediction_WORD_SLICES_BRANCH;
  reg        [1:0]    AlignerPlugin_logic_buffer_hm_Prediction_WORD_SLICES_TAKEN;
  reg        [38:0]   AlignerPlugin_logic_buffer_hm_Prediction_WORD_JUMP_PC;
  reg                 AlignerPlugin_logic_buffer_hm_Prediction_WORD_JUMPED;
  reg        [0:0]    AlignerPlugin_logic_buffer_hm_Prediction_WORD_JUMP_SLICE;
  wire       [63:0]   _zz_AlignerPlugin_logic_slices_data_0;
  wire                when_AlignerPlugin_l240;
  wire                when_AlignerPlugin_l241;
  wire                AlignerPlugin_logic_buffer_downFire;
  wire       [3:0]    AlignerPlugin_logic_buffer_usedMask;
  wire                AlignerPlugin_logic_buffer_haltUp;
  wire                when_AlignerPlugin_l256;
  wire       [1:0]    early0_EnvPlugin_logic_exe_privilege;
  wire       [1:0]    early0_EnvPlugin_logic_exe_xretPriv;
  reg                 early0_EnvPlugin_logic_exe_commit;
  wire                early0_EnvPlugin_logic_exe_retKo;
  wire                early0_EnvPlugin_logic_exe_vmaKo;
  wire                when_EnvPlugin_l86;
  wire                when_EnvPlugin_l95;
  wire                when_EnvPlugin_l110;
  wire                when_EnvPlugin_l119;
  wire                when_EnvPlugin_l123;
  reg                 PerformanceCounterPlugin_logic_readPort_valid;
  wire                PerformanceCounterPlugin_logic_readPort_ready;
  wire       [3:0]    PerformanceCounterPlugin_logic_readPort_address;
  wire       [63:0]   PerformanceCounterPlugin_logic_readPort_data;
  reg                 PerformanceCounterPlugin_logic_writePort_valid;
  wire                PerformanceCounterPlugin_logic_writePort_ready;
  wire       [3:0]    PerformanceCounterPlugin_logic_writePort_address;
  reg        [63:0]   PerformanceCounterPlugin_logic_writePort_data;
  wire                PmpPlugin_logic_isMachine;
  wire                PmpPlugin_logic_instructionShouldHit;
  wire                PmpPlugin_logic_dataShouldHit;
  wire                FetchL1Plugin_logic_pmpPort_logic_dataShouldHitPort;
  wire       [19:0]   FetchL1Plugin_logic_pmpPort_logic_torCmpAddress;
  wire                FetchL1Plugin_logic_pmpPort_logic_onEntries_0_instructionCheck;
  wire                FetchL1Plugin_logic_pmpPort_logic_onEntries_0_dataCheck;
  wire                FetchL1Plugin_logic_pmpPort_logic_onEntries_0_normalRwx;
  wire                FetchL1Plugin_logic_pmpPort_logic_onEntries_1_instructionCheck;
  wire                FetchL1Plugin_logic_pmpPort_logic_onEntries_1_dataCheck;
  wire                FetchL1Plugin_logic_pmpPort_logic_onEntries_1_normalRwx;
  wire                FetchL1Plugin_logic_pmpPort_logic_onEntries_2_instructionCheck;
  wire                FetchL1Plugin_logic_pmpPort_logic_onEntries_2_dataCheck;
  wire                FetchL1Plugin_logic_pmpPort_logic_onEntries_2_normalRwx;
  wire                FetchL1Plugin_logic_pmpPort_logic_onEntries_3_instructionCheck;
  wire                FetchL1Plugin_logic_pmpPort_logic_onEntries_3_dataCheck;
  wire                FetchL1Plugin_logic_pmpPort_logic_onEntries_3_normalRwx;
  wire       [3:0]    FetchL1Plugin_logic_pmpPort_logic_onCtrl_hits;
  wire       [3:0]    _zz_FetchL1Plugin_logic_pmpPort_logic_onCtrl_hits_bools_0;
  wire                FetchL1Plugin_logic_pmpPort_logic_onCtrl_hits_bools_0;
  wire                FetchL1Plugin_logic_pmpPort_logic_onCtrl_hits_bools_1;
  wire                FetchL1Plugin_logic_pmpPort_logic_onCtrl_hits_bools_2;
  wire                FetchL1Plugin_logic_pmpPort_logic_onCtrl_hits_bools_3;
  reg        [3:0]    _zz_FetchL1Plugin_logic_pmpPort_logic_onCtrl_oh;
  wire                FetchL1Plugin_logic_pmpPort_logic_onCtrl_hits_range_0_to_1;
  wire                FetchL1Plugin_logic_pmpPort_logic_onCtrl_hits_range_0_to_2;
  wire       [3:0]    FetchL1Plugin_logic_pmpPort_logic_onCtrl_oh;
  wire                _zz_fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_ACCESS_FAULT;
  wire                _zz_fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_ACCESS_FAULT_1;
  wire                _zz_fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_ACCESS_FAULT_2;
  wire                _zz_fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_ACCESS_FAULT_3;
  wire                LsuPlugin_logic_pmpPort_logic_dataShouldHitPort;
  wire       [19:0]   LsuPlugin_logic_pmpPort_logic_torCmpAddress;
  wire                LsuPlugin_logic_pmpPort_logic_onEntries_0_instructionCheck;
  wire                LsuPlugin_logic_pmpPort_logic_onEntries_0_dataCheck;
  wire                LsuPlugin_logic_pmpPort_logic_onEntries_0_normalRwx;
  wire                LsuPlugin_logic_pmpPort_logic_onEntries_1_instructionCheck;
  wire                LsuPlugin_logic_pmpPort_logic_onEntries_1_dataCheck;
  wire                LsuPlugin_logic_pmpPort_logic_onEntries_1_normalRwx;
  wire                LsuPlugin_logic_pmpPort_logic_onEntries_2_instructionCheck;
  wire                LsuPlugin_logic_pmpPort_logic_onEntries_2_dataCheck;
  wire                LsuPlugin_logic_pmpPort_logic_onEntries_2_normalRwx;
  wire                LsuPlugin_logic_pmpPort_logic_onEntries_3_instructionCheck;
  wire                LsuPlugin_logic_pmpPort_logic_onEntries_3_dataCheck;
  wire                LsuPlugin_logic_pmpPort_logic_onEntries_3_normalRwx;
  wire       [3:0]    LsuPlugin_logic_pmpPort_logic_onCtrl_hits;
  wire       [3:0]    _zz_LsuPlugin_logic_pmpPort_logic_onCtrl_hits_bools_0;
  wire                LsuPlugin_logic_pmpPort_logic_onCtrl_hits_bools_0;
  wire                LsuPlugin_logic_pmpPort_logic_onCtrl_hits_bools_1;
  wire                LsuPlugin_logic_pmpPort_logic_onCtrl_hits_bools_2;
  wire                LsuPlugin_logic_pmpPort_logic_onCtrl_hits_bools_3;
  reg        [3:0]    _zz_LsuPlugin_logic_pmpPort_logic_onCtrl_oh;
  wire                LsuPlugin_logic_pmpPort_logic_onCtrl_hits_range_0_to_1;
  wire                LsuPlugin_logic_pmpPort_logic_onCtrl_hits_range_0_to_2;
  wire       [3:0]    LsuPlugin_logic_pmpPort_logic_onCtrl_oh;
  wire                _zz_execute_ctrl4_down_LsuPlugin_logic_pmpPort_ACCESS_FAULT_lane0;
  wire                _zz_execute_ctrl4_down_LsuPlugin_logic_pmpPort_ACCESS_FAULT_lane0_1;
  wire                _zz_execute_ctrl4_down_LsuPlugin_logic_pmpPort_ACCESS_FAULT_lane0_2;
  wire                _zz_execute_ctrl4_down_LsuPlugin_logic_pmpPort_ACCESS_FAULT_lane0_3;
  wire                LsuCachelessAxi4Plugin_logic_bridge_down_arw_valid;
  wire                LsuCachelessAxi4Plugin_logic_bridge_down_arw_ready;
  wire       [31:0]   LsuCachelessAxi4Plugin_logic_bridge_down_arw_payload_addr;
  wire       [2:0]    LsuCachelessAxi4Plugin_logic_bridge_down_arw_payload_size;
  wire       [3:0]    LsuCachelessAxi4Plugin_logic_bridge_down_arw_payload_cache;
  wire       [2:0]    LsuCachelessAxi4Plugin_logic_bridge_down_arw_payload_prot;
  wire                LsuCachelessAxi4Plugin_logic_bridge_down_arw_payload_write;
  wire                LsuCachelessAxi4Plugin_logic_bridge_down_w_valid;
  wire                LsuCachelessAxi4Plugin_logic_bridge_down_w_ready;
  wire       [63:0]   LsuCachelessAxi4Plugin_logic_bridge_down_w_payload_data;
  wire       [7:0]    LsuCachelessAxi4Plugin_logic_bridge_down_w_payload_strb;
  wire                LsuCachelessAxi4Plugin_logic_bridge_down_w_payload_last;
  wire                LsuCachelessAxi4Plugin_logic_bridge_down_b_valid;
  reg                 LsuCachelessAxi4Plugin_logic_bridge_down_b_ready;
  wire       [1:0]    LsuCachelessAxi4Plugin_logic_bridge_down_b_payload_resp;
  wire                LsuCachelessAxi4Plugin_logic_bridge_down_r_valid;
  wire                LsuCachelessAxi4Plugin_logic_bridge_down_r_ready;
  wire       [63:0]   LsuCachelessAxi4Plugin_logic_bridge_down_r_payload_data;
  wire       [1:0]    LsuCachelessAxi4Plugin_logic_bridge_down_r_payload_resp;
  wire                LsuCachelessAxi4Plugin_logic_bridge_down_r_payload_last;
  wire                LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_valid;
  reg                 LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_ready;
  wire                LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_payload_write;
  wire       [31:0]   LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_payload_address;
  wire       [63:0]   LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_payload_data;
  wire       [1:0]    LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_payload_size;
  wire       [7:0]    LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_payload_mask;
  wire                LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_payload_io;
  wire                LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_payload_fromHart;
  wire       [15:0]   LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_payload_uopId;
  wire       [7:0]    LsuCachelessAxi4Plugin_logic_bridge_cmdHash;
  reg                 LsuCachelessAxi4Plugin_logic_bridge_tracker_pendings_0_valid;
  reg        [7:0]    LsuCachelessAxi4Plugin_logic_bridge_tracker_pendings_0_hash;
  reg        [7:0]    LsuCachelessAxi4Plugin_logic_bridge_tracker_pendings_0_mask;
  reg                 LsuCachelessAxi4Plugin_logic_bridge_tracker_pendings_0_io;
  wire                LsuCachelessAxi4Plugin_logic_bridge_tracker_pendings_0_hazard;
  wire                LsuCachelessAxi4Plugin_logic_bridge_tracker_hazard;
  wire                _zz_LsuPlugin_logic_bus_cmd_ready;
  wire                LsuPlugin_logic_bus_cmd_haltWhen_valid;
  wire                LsuPlugin_logic_bus_cmd_haltWhen_ready;
  wire                LsuPlugin_logic_bus_cmd_haltWhen_payload_write;
  wire       [31:0]   LsuPlugin_logic_bus_cmd_haltWhen_payload_address;
  wire       [63:0]   LsuPlugin_logic_bus_cmd_haltWhen_payload_data;
  wire       [1:0]    LsuPlugin_logic_bus_cmd_haltWhen_payload_size;
  wire       [7:0]    LsuPlugin_logic_bus_cmd_haltWhen_payload_mask;
  wire                LsuPlugin_logic_bus_cmd_haltWhen_payload_io;
  wire                LsuPlugin_logic_bus_cmd_haltWhen_payload_fromHart;
  wire       [15:0]   LsuPlugin_logic_bus_cmd_haltWhen_payload_uopId;
  wire                LsuCachelessAxi4Plugin_logic_bridge_cmdFork_valid;
  wire                LsuCachelessAxi4Plugin_logic_bridge_cmdFork_ready;
  wire                LsuCachelessAxi4Plugin_logic_bridge_cmdFork_payload_write;
  wire       [31:0]   LsuCachelessAxi4Plugin_logic_bridge_cmdFork_payload_address;
  wire       [63:0]   LsuCachelessAxi4Plugin_logic_bridge_cmdFork_payload_data;
  wire       [1:0]    LsuCachelessAxi4Plugin_logic_bridge_cmdFork_payload_size;
  wire       [7:0]    LsuCachelessAxi4Plugin_logic_bridge_cmdFork_payload_mask;
  wire                LsuCachelessAxi4Plugin_logic_bridge_cmdFork_payload_io;
  wire                LsuCachelessAxi4Plugin_logic_bridge_cmdFork_payload_fromHart;
  wire       [15:0]   LsuCachelessAxi4Plugin_logic_bridge_cmdFork_payload_uopId;
  wire                LsuCachelessAxi4Plugin_logic_bridge_dataFork_valid;
  reg                 LsuCachelessAxi4Plugin_logic_bridge_dataFork_ready;
  wire                LsuCachelessAxi4Plugin_logic_bridge_dataFork_payload_write;
  wire       [31:0]   LsuCachelessAxi4Plugin_logic_bridge_dataFork_payload_address;
  wire       [63:0]   LsuCachelessAxi4Plugin_logic_bridge_dataFork_payload_data;
  wire       [1:0]    LsuCachelessAxi4Plugin_logic_bridge_dataFork_payload_size;
  wire       [7:0]    LsuCachelessAxi4Plugin_logic_bridge_dataFork_payload_mask;
  wire                LsuCachelessAxi4Plugin_logic_bridge_dataFork_payload_io;
  wire                LsuCachelessAxi4Plugin_logic_bridge_dataFork_payload_fromHart;
  wire       [15:0]   LsuCachelessAxi4Plugin_logic_bridge_dataFork_payload_uopId;
  reg                 LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_fork2_logic_linkEnable_0;
  reg                 LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_fork2_logic_linkEnable_1;
  wire                when_Stream_l1253_2;
  wire                when_Stream_l1253_3;
  wire                LsuCachelessAxi4Plugin_logic_bridge_cmdFork_fire;
  wire                LsuCachelessAxi4Plugin_logic_bridge_dataFork_fire;
  wire                when_Stream_l581_1;
  reg                 LsuCachelessAxi4Plugin_logic_bridge_dataStage_valid;
  wire                LsuCachelessAxi4Plugin_logic_bridge_dataStage_ready;
  wire                LsuCachelessAxi4Plugin_logic_bridge_dataStage_payload_write;
  wire       [31:0]   LsuCachelessAxi4Plugin_logic_bridge_dataStage_payload_address;
  wire       [63:0]   LsuCachelessAxi4Plugin_logic_bridge_dataStage_payload_data;
  wire       [1:0]    LsuCachelessAxi4Plugin_logic_bridge_dataStage_payload_size;
  wire       [7:0]    LsuCachelessAxi4Plugin_logic_bridge_dataStage_payload_mask;
  wire                LsuCachelessAxi4Plugin_logic_bridge_dataStage_payload_io;
  wire                LsuCachelessAxi4Plugin_logic_bridge_dataStage_payload_fromHart;
  wire       [15:0]   LsuCachelessAxi4Plugin_logic_bridge_dataStage_payload_uopId;
  wire       [31:0]   LsuPlugin_pmaBuilder_l1_addressBits;
  wire       [0:0]    LsuPlugin_pmaBuilder_l1_argsBits;
  wire                _zz_LsuPlugin_logic_onPma_cached_rsp_io;
  wire                LsuPlugin_pmaBuilder_l1_onTransfers_0_addressHit;
  wire                LsuPlugin_pmaBuilder_l1_onTransfers_0_argsHit;
  wire                LsuPlugin_pmaBuilder_l1_onTransfers_0_hit;
  wire       [31:0]   LsuPlugin_pmaBuilder_io_addressBits;
  wire       [2:0]    LsuPlugin_pmaBuilder_io_argsBits;
  wire                LsuPlugin_pmaBuilder_io_onTransfers_0_addressHit;
  wire                LsuPlugin_pmaBuilder_io_onTransfers_0_argsHit;
  wire                LsuPlugin_pmaBuilder_io_onTransfers_0_hit;
  wire                CsrRamPlugin_setup_initPort_valid;
  wire                CsrRamPlugin_setup_initPort_ready;
  wire       [3:0]    CsrRamPlugin_setup_initPort_address;
  wire       [63:0]   CsrRamPlugin_setup_initPort_data;
  wire                early0_BranchPlugin_logic_alu_expectedMsb;
  wire       [24:0]   _zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0;
  wire       [2:0]    switch_Misc_l245_1;
  reg                 _zz_execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0;
  reg                 _zz_execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0_1;
  wire                early0_BranchPlugin_logic_jumpLogic_wrongCond;
  wire                early0_BranchPlugin_logic_jumpLogic_needFix;
  wire                early0_BranchPlugin_logic_jumpLogic_doIt;
  wire       [11:0]   early0_BranchPlugin_logic_jumpLogic_history_fetched;
  wire       [11:0]   early0_BranchPlugin_logic_jumpLogic_history_next;
  wire       [0:0]    early0_BranchPlugin_logic_jumpLogic_history_slice;
  wire       [11:0]   early0_BranchPlugin_logic_jumpLogic_history_shifter;
  wire                when_BranchPlugin_l213;
  wire                when_BranchPlugin_l218;
  wire                early0_BranchPlugin_logic_jumpLogic_rdLink;
  wire                early0_BranchPlugin_logic_jumpLogic_rs1Link;
  wire                early0_BranchPlugin_logic_jumpLogic_rdEquRs1;
  wire                early0_BranchPlugin_logic_jumpLogic_learn_valid;
  wire                early0_BranchPlugin_logic_jumpLogic_learn_ready;
  wire       [38:0]   early0_BranchPlugin_logic_jumpLogic_learn_payload_pcOnLastSlice;
  wire       [38:0]   early0_BranchPlugin_logic_jumpLogic_learn_payload_pcTarget;
  wire                early0_BranchPlugin_logic_jumpLogic_learn_payload_taken;
  wire                early0_BranchPlugin_logic_jumpLogic_learn_payload_isBranch;
  wire                early0_BranchPlugin_logic_jumpLogic_learn_payload_isPush;
  wire                early0_BranchPlugin_logic_jumpLogic_learn_payload_isPop;
  wire                early0_BranchPlugin_logic_jumpLogic_learn_payload_wasWrong;
  wire                early0_BranchPlugin_logic_jumpLogic_learn_payload_badPredictedTarget;
  wire       [11:0]   early0_BranchPlugin_logic_jumpLogic_learn_payload_history;
  wire       [15:0]   early0_BranchPlugin_logic_jumpLogic_learn_payload_uopId;
  wire       [1:0]    early0_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    early0_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  wire                CsrRamPlugin_csrMapper_read_valid;
  wire                CsrRamPlugin_csrMapper_read_ready;
  wire       [3:0]    CsrRamPlugin_csrMapper_read_address;
  wire       [63:0]   CsrRamPlugin_csrMapper_read_data;
  wire                CsrRamPlugin_csrMapper_write_valid;
  wire                CsrRamPlugin_csrMapper_write_ready;
  wire       [3:0]    CsrRamPlugin_csrMapper_write_address;
  wire       [63:0]   CsrRamPlugin_csrMapper_write_data;
  wire                LearnPlugin_logic_learn_valid;
  wire       [38:0]   LearnPlugin_logic_learn_payload_pcOnLastSlice;
  wire       [38:0]   LearnPlugin_logic_learn_payload_pcTarget;
  wire                LearnPlugin_logic_learn_payload_taken;
  wire                LearnPlugin_logic_learn_payload_isBranch;
  wire                LearnPlugin_logic_learn_payload_isPush;
  wire                LearnPlugin_logic_learn_payload_isPop;
  wire                LearnPlugin_logic_learn_payload_wasWrong;
  wire                LearnPlugin_logic_learn_payload_badPredictedTarget;
  wire       [11:0]   LearnPlugin_logic_learn_payload_history;
  wire       [15:0]   LearnPlugin_logic_learn_payload_uopId;
  wire       [1:0]    LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  wire                LearnPlugin_logic_buffered_0_valid;
  wire                LearnPlugin_logic_buffered_0_ready;
  wire       [38:0]   LearnPlugin_logic_buffered_0_payload_pcOnLastSlice;
  wire       [38:0]   LearnPlugin_logic_buffered_0_payload_pcTarget;
  wire                LearnPlugin_logic_buffered_0_payload_taken;
  wire                LearnPlugin_logic_buffered_0_payload_isBranch;
  wire                LearnPlugin_logic_buffered_0_payload_isPush;
  wire                LearnPlugin_logic_buffered_0_payload_isPop;
  wire                LearnPlugin_logic_buffered_0_payload_wasWrong;
  wire                LearnPlugin_logic_buffered_0_payload_badPredictedTarget;
  wire       [11:0]   LearnPlugin_logic_buffered_0_payload_history;
  wire       [15:0]   LearnPlugin_logic_buffered_0_payload_uopId;
  wire       [1:0]    LearnPlugin_logic_buffered_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    LearnPlugin_logic_buffered_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  wire                LearnPlugin_logic_arbitrated_valid;
  wire                LearnPlugin_logic_arbitrated_ready;
  wire       [38:0]   LearnPlugin_logic_arbitrated_payload_pcOnLastSlice;
  wire       [38:0]   LearnPlugin_logic_arbitrated_payload_pcTarget;
  wire                LearnPlugin_logic_arbitrated_payload_taken;
  wire                LearnPlugin_logic_arbitrated_payload_isBranch;
  wire                LearnPlugin_logic_arbitrated_payload_isPush;
  wire                LearnPlugin_logic_arbitrated_payload_isPop;
  wire                LearnPlugin_logic_arbitrated_payload_wasWrong;
  wire                LearnPlugin_logic_arbitrated_payload_badPredictedTarget;
  wire       [11:0]   LearnPlugin_logic_arbitrated_payload_history;
  wire       [15:0]   LearnPlugin_logic_arbitrated_payload_uopId;
  wire       [1:0]    LearnPlugin_logic_arbitrated_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    LearnPlugin_logic_arbitrated_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  wire                LearnPlugin_logic_arbitrated_toFlow_valid;
  wire       [38:0]   LearnPlugin_logic_arbitrated_toFlow_payload_pcOnLastSlice;
  wire       [38:0]   LearnPlugin_logic_arbitrated_toFlow_payload_pcTarget;
  wire                LearnPlugin_logic_arbitrated_toFlow_payload_taken;
  wire                LearnPlugin_logic_arbitrated_toFlow_payload_isBranch;
  wire                LearnPlugin_logic_arbitrated_toFlow_payload_isPush;
  wire                LearnPlugin_logic_arbitrated_toFlow_payload_isPop;
  wire                LearnPlugin_logic_arbitrated_toFlow_payload_wasWrong;
  wire                LearnPlugin_logic_arbitrated_toFlow_payload_badPredictedTarget;
  wire       [11:0]   LearnPlugin_logic_arbitrated_toFlow_payload_history;
  wire       [15:0]   LearnPlugin_logic_arbitrated_toFlow_payload_uopId;
  wire       [1:0]    LearnPlugin_logic_arbitrated_toFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    LearnPlugin_logic_arbitrated_toFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  reg        [15:0]   DecoderPlugin_logic_harts_0_uopId;
  wire                when_DecoderPlugin_l143;
  wire       [0:0]    DecoderPlugin_logic_interrupt_async;
  wire                when_DecoderPlugin_l151;
  reg        [0:0]    DecoderPlugin_logic_interrupt_buffered;
  wire                when_DecoderPlugin_l187;
  wire                when_DecoderPlugin_l187_1;
  wire                DecoderPlugin_logic_laneLogic_0_interruptPending;
  reg                 DecoderPlugin_logic_laneLogic_0_trapPort_valid;
  reg                 DecoderPlugin_logic_laneLogic_0_trapPort_payload_exception;
  wire       [38:0]   DecoderPlugin_logic_laneLogic_0_trapPort_payload_tval;
  reg        [3:0]    DecoderPlugin_logic_laneLogic_0_trapPort_payload_code;
  wire       [2:0]    DecoderPlugin_logic_laneLogic_0_trapPort_payload_arg;
  wire       [0:0]    DecoderPlugin_logic_laneLogic_0_trapPort_payload_laneAge;
  wire                DecoderPlugin_logic_laneLogic_0_fixer_isJb;
  wire                DecoderPlugin_logic_laneLogic_0_fixer_doIt;
  wire                DecoderPlugin_logic_laneLogic_0_completionPort_valid;
  wire       [15:0]   DecoderPlugin_logic_laneLogic_0_completionPort_payload_uopId;
  wire                DecoderPlugin_logic_laneLogic_0_completionPort_payload_trap;
  wire                DecoderPlugin_logic_laneLogic_0_completionPort_payload_commit;
  reg                 decode_ctrls_1_up_LANE_SEL_0_regNext;
  wire                when_CtrlLaneApi_l50_1;
  wire                when_DecoderPlugin_l229;
  wire                DecoderPlugin_logic_laneLogic_0_flushPort_valid;
  wire       [15:0]   DecoderPlugin_logic_laneLogic_0_flushPort_payload_uopId;
  wire                DecoderPlugin_logic_laneLogic_0_flushPort_payload_self;
  wire                when_DecoderPlugin_l247;
  wire       [15:0]   DecoderPlugin_logic_laneLogic_0_uopIdBase;
  wire                DispatchPlugin_logic_candidates_0_ctx_valid;
  reg        [0:0]    DispatchPlugin_logic_candidates_0_ctx_laneLayerHits;
  wire       [31:0]   DispatchPlugin_logic_candidates_0_ctx_uop;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_JUMPED;
  wire       [38:0]   DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_JUMPED_PC;
  wire       [1:0]    DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_SLICES_TAKEN;
  wire       [1:0]    DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_SLICES_BRANCH;
  wire       [1:0]    DispatchPlugin_logic_candidates_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    DispatchPlugin_logic_candidates_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_1;
  wire       [11:0]   DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_BRANCH_HISTORY;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_FENCE_OLDER;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_MAY_FLUSH;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_DONT_FLUSH;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES;
  wire       [0:0]    DispatchPlugin_logic_candidates_0_ctx_hm_Decode_INSTRUCTION_SLICE_COUNT;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_3;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_4;
  wire       [38:0]   DispatchPlugin_logic_candidates_0_ctx_hm_PC;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_TRAP;
  wire       [15:0]   DispatchPlugin_logic_candidates_0_ctx_hm_Decode_UOP_ID;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_RS1_ENABLE;
  wire       [4:0]    DispatchPlugin_logic_candidates_0_ctx_hm_RS1_PHYS;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_RS2_ENABLE;
  wire       [4:0]    DispatchPlugin_logic_candidates_0_ctx_hm_RS2_PHYS;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_RD_ENABLE;
  wire       [4:0]    DispatchPlugin_logic_candidates_0_ctx_hm_RD_PHYS;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_0_fire;
  wire                DispatchPlugin_logic_candidates_0_cancel;
  wire       [0:0]    DispatchPlugin_logic_candidates_0_rsHazards;
  wire       [0:0]    DispatchPlugin_logic_candidates_0_reservationHazards;
  wire                DispatchPlugin_logic_candidates_0_flushHazards;
  wire                DispatchPlugin_logic_candidates_0_fenceOlderHazards;
  wire                DispatchPlugin_logic_candidates_0_moving;
  wire                DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard;
  wire                DispatchPlugin_logic_reservationChecker_0_onLl_0_hit;
  wire                DispatchPlugin_logic_flushChecker_0_executeCheck_0_hits_0;
  wire                DispatchPlugin_logic_flushChecker_0_executeCheck_0_hits_1;
  wire                DispatchPlugin_logic_flushChecker_0_oldersHazard;
  wire       [0:0]    DispatchPlugin_logic_fenceChecker_olderInflights;
  wire                DispatchPlugin_logic_feeds_0_sending;
  reg                 DispatchPlugin_logic_feeds_0_sent;
  wire                when_DispatchPlugin_l368;
  wire       [0:0]    DispatchPlugin_logic_scheduler_eusFree_0;
  wire       [0:0]    DispatchPlugin_logic_scheduler_eusFree_1;
  wire       [0:0]    DispatchPlugin_logic_scheduler_hartFree_0;
  wire       [0:0]    DispatchPlugin_logic_scheduler_hartFree_1;
  wire                DispatchPlugin_logic_scheduler_arbiters_0_candHazard;
  wire       [0:0]    DispatchPlugin_logic_scheduler_arbiters_0_layersHits;
  wire                DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_0;
  wire       [0:0]    _zz_DispatchPlugin_logic_scheduler_arbiters_0_layerOh;
  wire       [0:0]    DispatchPlugin_logic_scheduler_arbiters_0_layerOh;
  wire       [0:0]    DispatchPlugin_logic_scheduler_arbiters_0_eusOh;
  wire                DispatchPlugin_logic_scheduler_arbiters_0_doIt;
  wire       [0:0]    DispatchPlugin_logic_inserter_0_oh;
  wire                DispatchPlugin_logic_inserter_0_trap;
  wire                when_DispatchPlugin_l439;
  wire       [0:0]    DispatchPlugin_logic_inserter_0_layerOhUnfiltred;
  wire                DispatchPlugin_logic_inserter_0_layer_0_1;
  wire                DispatchPlugin_logic_events_frontendStall;
  wire                DispatchPlugin_logic_events_backendStall;
  wire       [3:0]    CsrRamPlugin_csrMapper_ramAddress;
  wire       [11:0]   _zz_CsrRamPlugin_csrMapper_ramAddress;
  reg                 CsrRamPlugin_csrMapper_withRead;
  wire                when_CsrRamPlugin_l90;
  reg                 CsrRamPlugin_csrMapper_doWrite;
  reg                 CsrRamPlugin_csrMapper_fired;
  wire                when_CsrRamPlugin_l97;
  wire                when_CsrRamPlugin_l101;
  wire       [12:0]   _zz_GSharePlugin_logic_onLearn_hash;
  wire       [12:0]   GSharePlugin_logic_onLearn_hash;
  wire       [1:0]    GSharePlugin_logic_onLearn_updated_0;
  wire       [1:0]    GSharePlugin_logic_onLearn_updated_1;
  wire       [1:0]    GSharePlugin_logic_onLearn_incrValue;
  reg                 GSharePlugin_logic_onLearn_overflow;
  wire                when_GSharePlugin_l119;
  wire                when_GSharePlugin_l119_1;
  wire       [15:0]   BtbPlugin_logic_onLearn_hash;
  wire       [1:0]    lane0_integer_WriteBackPlugin_logic_stages_0_hits;
  wire       [63:0]   lane0_integer_WriteBackPlugin_logic_stages_0_muxed;
  wire                lane0_integer_WriteBackPlugin_logic_stages_0_write_valid;
  wire       [15:0]   lane0_integer_WriteBackPlugin_logic_stages_0_write_payload_uopId;
  wire       [63:0]   lane0_integer_WriteBackPlugin_logic_stages_0_write_payload_data;
  wire       [0:0]    lane0_integer_WriteBackPlugin_logic_stages_1_hits;
  wire       [63:0]   lane0_integer_WriteBackPlugin_logic_stages_1_muxed;
  wire       [63:0]   lane0_integer_WriteBackPlugin_logic_stages_1_merged;
  wire                lane0_integer_WriteBackPlugin_logic_stages_1_write_valid;
  wire       [15:0]   lane0_integer_WriteBackPlugin_logic_stages_1_write_payload_uopId;
  wire       [63:0]   lane0_integer_WriteBackPlugin_logic_stages_1_write_payload_data;
  wire       [0:0]    lane0_integer_WriteBackPlugin_logic_stages_2_hits;
  wire       [63:0]   lane0_integer_WriteBackPlugin_logic_stages_2_muxed;
  wire       [63:0]   lane0_integer_WriteBackPlugin_logic_stages_2_merged;
  wire                lane0_integer_WriteBackPlugin_logic_stages_2_write_valid;
  wire       [15:0]   lane0_integer_WriteBackPlugin_logic_stages_2_write_payload_uopId;
  wire       [63:0]   lane0_integer_WriteBackPlugin_logic_stages_2_write_payload_data;
  wire                lane0_integer_WriteBackPlugin_logic_write_port_valid;
  wire       [4:0]    lane0_integer_WriteBackPlugin_logic_write_port_address;
  wire       [63:0]   lane0_integer_WriteBackPlugin_logic_write_port_data;
  wire       [15:0]   lane0_integer_WriteBackPlugin_logic_write_port_uopId;
  wire                _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0;
  wire                _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0;
  wire                _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_1;
  wire                TrapPlugin_logic_initHold;
  reg                 decode_ctrls_1_up_LANE_SEL_0_regNext_1;
  wire                when_CtrlLaneApi_l50_2;
  wire                WhiteboxerPlugin_logic_serializeds_0_fire;
  wire       [9:0]    WhiteboxerPlugin_logic_serializeds_0_decodeId;
  wire       [15:0]   WhiteboxerPlugin_logic_serializeds_0_microOpId;
  wire       [31:0]   WhiteboxerPlugin_logic_serializeds_0_microOp;
  reg                 execute_ctrl0_down_LANE_SEL_lane0_regNext;
  wire                when_CtrlLaneApi_l50_3;
  wire                WhiteboxerPlugin_logic_dispatches_0_fire;
  wire       [15:0]   WhiteboxerPlugin_logic_dispatches_0_microOpId;
  reg                 execute_ctrl2_down_LANE_SEL_lane0_regNext;
  wire                when_CtrlLaneApi_l50_4;
  wire                WhiteboxerPlugin_logic_executes_0_fire;
  wire       [15:0]   WhiteboxerPlugin_logic_executes_0_microOpId;
  wire                WhiteboxerPlugin_logic_csr_access_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_csr_access_payload_uopId;
  wire       [11:0]   WhiteboxerPlugin_logic_csr_access_payload_address;
  wire       [63:0]   WhiteboxerPlugin_logic_csr_access_payload_write;
  wire       [63:0]   WhiteboxerPlugin_logic_csr_access_payload_read;
  wire                WhiteboxerPlugin_logic_csr_access_payload_writeDone;
  wire                WhiteboxerPlugin_logic_csr_access_payload_readDone;
  wire       [15:0]   BtbPlugin_logic_onForget_hash;
  wire                fetch_logic_ctrls_0_haltRequest_BtbPlugin_l200;
  wire       [1:0]    BtbPlugin_logic_predictions;
  wire       [0:0]    BtbPlugin_logic_applyIt_chunksMask;
  wire       [0:0]    BtbPlugin_logic_applyIt_chunksTakenOh;
  wire                BtbPlugin_logic_applyIt_needIt;
  reg                 BtbPlugin_logic_applyIt_correctionSent;
  wire                when_BtbPlugin_l233;
  wire                BtbPlugin_logic_applyIt_doIt;
  wire       [15:0]   BtbPlugin_logic_applyIt_entry_hash;
  wire       [0:0]    BtbPlugin_logic_applyIt_entry_sliceLow;
  wire       [37:0]   BtbPlugin_logic_applyIt_entry_pcTarget;
  wire                BtbPlugin_logic_applyIt_entry_isBranch;
  wire                BtbPlugin_logic_applyIt_entry_isPush;
  wire                BtbPlugin_logic_applyIt_entry_isPop;
  reg        [37:0]   BtbPlugin_logic_applyIt_pcTarget;
  wire       [0:0]    BtbPlugin_logic_applyIt_doItSlice;
  wire                BtbPlugin_logic_applyIt_rasLogic_pushValid;
  reg        [38:0]   BtbPlugin_logic_applyIt_rasLogic_pushPc;
  wire                when_BtbPlugin_l246;
  wire       [11:0]   BtbPlugin_logic_applyIt_history_layers_0_history;
  wire                BtbPlugin_logic_applyIt_history_layers_0_valid;
  wire       [11:0]   BtbPlugin_logic_applyIt_history_layers_1_history;
  wire                BtbPlugin_logic_applyIt_history_layers_1_valid;
  wire                BtbPlugin_logic_applyIt_history_layersLogic_0_doIt;
  wire       [11:0]   BtbPlugin_logic_applyIt_history_layersLogic_0_shifted;
  reg                 TrapPlugin_logic_harts_0_crsPorts_read_valid;
  wire                TrapPlugin_logic_harts_0_crsPorts_read_ready;
  reg        [3:0]    TrapPlugin_logic_harts_0_crsPorts_read_address;
  wire       [63:0]   TrapPlugin_logic_harts_0_crsPorts_read_data;
  wire                AlignerPlugin_logic_buffer_flushIt;
  wire                AlignerPlugin_logic_buffer_readers_0_firstFromBuffer;
  wire                AlignerPlugin_logic_buffer_readers_0_lastFromBuffer;
  wire       [3:0]    _zz_AlignerPlugin_logic_extractors_0_ctx_instruction;
  wire                _zz_AlignerPlugin_logic_extractors_0_ctx_pc;
  wire                decode_logic_flushes_0_onLanes_0_doIt;
  wire                decode_logic_flushes_1_onLanes_0_doIt;
  reg                 TrapPlugin_logic_harts_0_crsPorts_write_valid;
  wire                TrapPlugin_logic_harts_0_crsPorts_write_ready;
  reg        [3:0]    TrapPlugin_logic_harts_0_crsPorts_write_address;
  reg        [63:0]   TrapPlugin_logic_harts_0_crsPorts_write_data;
  wire       [3:0]    TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_0_id;
  wire       [3:0]    TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_0_priority;
  wire       [1:0]    TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_0_privilege;
  wire                TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_0_valid;
  wire       [3:0]    TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_1_id;
  wire       [3:0]    TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_1_priority;
  wire       [1:0]    TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_1_privilege;
  wire                TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_1_valid;
  wire       [3:0]    TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_2_id;
  wire       [3:0]    TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_2_priority;
  wire       [1:0]    TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_2_privilege;
  wire                TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_2_valid;
  wire                _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_triggered_id;
  wire       [3:0]    _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_triggered_priority;
  wire       [1:0]    _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_triggered_privilege;
  wire                _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_triggered_valid;
  wire                _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_triggered_id_1;
  reg        [3:0]    TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_triggered_id;
  reg        [3:0]    TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_triggered_priority;
  reg        [1:0]    TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_triggered_privilege;
  reg                 TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_triggered_valid;
  wire       [3:0]    TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_0_id;
  wire       [3:0]    TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_0_priority;
  wire       [1:0]    TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_0_privilege;
  wire                TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_0_valid;
  wire       [3:0]    TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_1_id;
  wire       [3:0]    TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_1_priority;
  wire       [1:0]    TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_1_privilege;
  wire                TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_1_valid;
  wire       [3:0]    TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_2_id;
  wire       [3:0]    TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_2_priority;
  wire       [1:0]    TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_2_privilege;
  wire                TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_2_valid;
  wire       [3:0]    TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_3_id;
  wire       [3:0]    TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_3_priority;
  wire       [1:0]    TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_3_privilege;
  wire                TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_3_valid;
  wire       [3:0]    TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_4_id;
  wire       [3:0]    TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_4_priority;
  wire       [1:0]    TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_4_privilege;
  wire                TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_4_valid;
  wire       [3:0]    TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_5_id;
  wire       [3:0]    TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_5_priority;
  wire       [1:0]    TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_5_privilege;
  wire                TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_5_valid;
  wire                _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id;
  wire       [3:0]    _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_1;
  wire       [1:0]    _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_2;
  wire                _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_3;
  wire                _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_4;
  wire       [3:0]    _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_5;
  wire       [1:0]    _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_6;
  wire                _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_7;
  wire                _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_8;
  wire       [3:0]    _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_priority;
  wire       [1:0]    _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_privilege;
  wire                _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_valid;
  wire                _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_9;
  wire       [3:0]    _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_priority_1;
  wire       [1:0]    _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_privilege_1;
  wire                _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_valid_1;
  wire                _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_10;
  reg        [3:0]    TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id;
  reg        [3:0]    TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_priority;
  reg        [1:0]    TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_privilege;
  reg                 TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_valid;
  wire       [3:0]    TrapPlugin_logic_harts_0_interrupt_xtopi_0_int;
  wire       [3:0]    TrapPlugin_logic_harts_0_interrupt_xtopi_1_int;
  wire       [1:0]    _zz_TrapPlugin_logic_harts_0_interrupt_result_privilege;
  wire                _zz_TrapPlugin_logic_harts_0_interrupt_result_valid;
  wire       [1:0]    _zz_TrapPlugin_logic_harts_0_interrupt_result_privilege_1;
  wire                _zz_TrapPlugin_logic_harts_0_interrupt_result_valid_1;
  wire                _zz_TrapPlugin_logic_harts_0_interrupt_result_id;
  wire       [3:0]    TrapPlugin_logic_harts_0_interrupt_result_id;
  wire       [3:0]    TrapPlugin_logic_harts_0_interrupt_result_priority;
  wire       [1:0]    TrapPlugin_logic_harts_0_interrupt_result_privilege;
  wire                TrapPlugin_logic_harts_0_interrupt_result_valid;
  wire                TrapPlugin_logic_harts_0_interrupt_valid;
  wire       [3:0]    TrapPlugin_logic_harts_0_interrupt_code;
  wire       [1:0]    TrapPlugin_logic_harts_0_interrupt_targetPrivilege;
  reg                 TrapPlugin_logic_harts_0_interrupt_validBuffer;
  wire                TrapPlugin_logic_harts_0_interrupt_pendingInterrupt;
  wire                when_TrapPlugin_l269;
  wire                _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid;
  wire                _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_valid;
  wire                _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_valid;
  wire                _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid_1;
  wire                _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid;
  wire                TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_valid;
  wire                TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_exception;
  wire       [38:0]   TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_tval;
  wire       [3:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_code;
  wire       [2:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_arg;
  wire                TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid;
  wire                TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_exception;
  wire       [38:0]   TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_tval;
  wire       [3:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_code;
  wire       [2:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_arg;
  wire       [1:0]    _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_exception;
  wire       [46:0]   _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_exception_1;
  wire                TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid;
  wire                TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_exception;
  wire       [38:0]   TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_tval;
  wire       [3:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_code;
  wire       [2:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_arg;
  wire                TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_valid;
  wire                TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_exception;
  wire       [38:0]   TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_tval;
  wire       [3:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_code;
  wire       [2:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_arg;
  wire       [3:0]    _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh;
  wire                _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_1;
  wire                _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_2;
  wire                _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_3;
  reg        [3:0]    _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_4;
  wire       [3:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_oh;
  wire                TrapPlugin_logic_harts_0_trap_pending_arbiter_down_valid;
  wire                TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception;
  wire       [38:0]   TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_tval;
  wire       [3:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_code;
  wire       [2:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_arg;
  wire       [46:0]   _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception;
  reg                 TrapPlugin_logic_harts_0_trap_pending_state_exception;
  reg        [38:0]   TrapPlugin_logic_harts_0_trap_pending_state_tval;
  reg        [3:0]    TrapPlugin_logic_harts_0_trap_pending_state_code;
  reg        [2:0]    TrapPlugin_logic_harts_0_trap_pending_state_arg;
  reg        [38:0]   TrapPlugin_logic_harts_0_trap_pending_pc;
  reg        [11:0]   TrapPlugin_logic_harts_0_trap_pending_history;
  reg        [1:0]    TrapPlugin_logic_harts_0_trap_pending_slices;
  wire       [1:0]    TrapPlugin_logic_harts_0_trap_pending_xret_sourcePrivilege;
  reg        [1:0]    TrapPlugin_logic_harts_0_trap_pending_xret_targetPrivilege;
  reg        [1:0]    TrapPlugin_logic_harts_0_trap_exception_exceptionTargetPrivilegeUncapped;
  wire       [3:0]    TrapPlugin_logic_harts_0_trap_exception_code;
  wire                when_TrapPlugin_l306;
  wire                when_TrapPlugin_l306_1;
  wire                when_TrapPlugin_l306_2;
  wire                when_TrapPlugin_l306_3;
  wire                when_TrapPlugin_l306_4;
  wire                when_TrapPlugin_l306_5;
  wire                when_TrapPlugin_l306_6;
  wire       [1:0]    TrapPlugin_logic_harts_0_trap_exception_targetPrivilege;
  wire                execute_lane0_ctrls_5_upIsCancel;
  wire                execute_lane0_ctrls_5_downIsCancel;
  wire       [0:0]    TrapPlugin_logic_harts_0_trap_trigger_oh;
  wire                TrapPlugin_logic_harts_0_trap_trigger_valid;
  reg                 TrapPlugin_logic_harts_0_trap_whitebox_trap;
  reg                 TrapPlugin_logic_harts_0_trap_whitebox_interrupt;
  reg        [3:0]    TrapPlugin_logic_harts_0_trap_whitebox_code;
  reg                 TrapPlugin_logic_harts_0_trap_historyPort_valid;
  wire       [11:0]   TrapPlugin_logic_harts_0_trap_historyPort_payload_history;
  reg                 TrapPlugin_logic_harts_0_trap_pcPort_valid;
  wire                TrapPlugin_logic_harts_0_trap_pcPort_payload_fault;
  reg        [38:0]   TrapPlugin_logic_harts_0_trap_pcPort_payload_pc;
  wire                PcPlugin_logic_harts_0_aggregator_sortedByPriority_0_laneValid;
  wire                TrapPlugin_logic_harts_0_trap_fsm_wantExit;
  reg                 TrapPlugin_logic_harts_0_trap_fsm_wantStart;
  wire                TrapPlugin_logic_harts_0_trap_fsm_wantKill;
  wire                TrapPlugin_logic_harts_0_trap_fsm_inflightTrap;
  wire                TrapPlugin_logic_harts_0_trap_fsm_holdPort;
  reg                 TrapPlugin_logic_harts_0_trap_fsm_wfi;
  reg                 TrapPlugin_logic_harts_0_trap_fsm_buffer_sampleIt;
  reg                 TrapPlugin_logic_harts_0_trap_fsm_buffer_i_valid;
  reg        [3:0]    TrapPlugin_logic_harts_0_trap_fsm_buffer_i_code;
  reg        [1:0]    TrapPlugin_logic_harts_0_trap_fsm_buffer_i_targetPrivilege;
  wire                TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_interrupt;
  wire       [1:0]    TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_targetPrivilege;
  wire       [38:0]   TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_tval;
  wire       [3:0]    TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_code;
  wire                TrapPlugin_logic_harts_0_trap_fsm_resetToRunConditions_0;
  reg                 TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_cmd_valid;
  wire                TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_cmd_ready;
  wire       [38:0]   bits_address;
  wire       [0:0]    bits_storageId;
  wire                bits_storageEnable;
  reg                 TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_valid;
  reg                 bits_pageFault;
  reg                 bits_accessFault;
  reg                 bits_ae_ptw;
  reg                 bits_ae_final;
  reg                 bits_pf;
  wire                bits_gf;
  wire                bits_hr;
  wire                bits_hw;
  wire                bits_hx;
  wire       [19:0]   bits_pte_ppn;
  wire                bits_pte_d;
  wire                bits_pte_a;
  wire                bits_pte_g;
  wire                bits_pte_u;
  wire                bits_pte_x;
  wire                bits_pte_w;
  wire                bits_pte_r;
  wire                bits_pte_v;
  reg        [1:0]    bits_level;
  reg                 TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidate_cmd_valid;
  wire                TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidate_cmd_ready;
  reg                 TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidated;
  wire                TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidate_cmd_fire;
  wire                when_TrapPlugin_l399;
  reg        [38:0]   TrapPlugin_logic_harts_0_trap_fsm_jumpTarget;
  wire       [1:0]    TrapPlugin_logic_harts_0_trap_fsm_jumpOffset;
  reg                 TrapPlugin_logic_harts_0_trap_fsm_trapEnterDebug;
  wire                TrapPlugin_logic_harts_0_trap_fsm_triggerEbreak;
  reg                 TrapPlugin_logic_harts_0_trap_fsm_triggerEbreakReg;
  wire                when_TrapPlugin_l602;
  reg        [63:0]   TrapPlugin_logic_harts_0_trap_fsm_readed;
  wire       [1:0]    TrapPlugin_logic_harts_0_trap_fsm_xretPrivilege;
  wire                PcPlugin_logic_forcedSpawn;
  reg        [9:0]    PcPlugin_logic_harts_0_self_id;
  wire                PcPlugin_logic_harts_0_self_flow_valid;
  wire                PcPlugin_logic_harts_0_self_flow_payload_fault;
  wire       [38:0]   PcPlugin_logic_harts_0_self_flow_payload_pc;
  wire                PcPlugin_logic_harts_0_aggregator_sortedByPriority_3_laneValid;
  reg                 PcPlugin_logic_harts_0_self_increment;
  reg                 PcPlugin_logic_harts_0_self_fault;
  reg        [38:0]   PcPlugin_logic_harts_0_self_state;
  wire       [38:0]   PcPlugin_logic_harts_0_self_pc;
  wire                PcPlugin_logic_harts_0_aggregator_valids_0;
  wire                PcPlugin_logic_harts_0_aggregator_valids_1;
  wire                PcPlugin_logic_harts_0_aggregator_valids_2;
  wire                PcPlugin_logic_harts_0_aggregator_valids_3;
  wire       [3:0]    _zz_PcPlugin_logic_harts_0_aggregator_oh;
  wire                _zz_PcPlugin_logic_harts_0_aggregator_oh_1;
  wire                _zz_PcPlugin_logic_harts_0_aggregator_oh_2;
  wire                _zz_PcPlugin_logic_harts_0_aggregator_oh_3;
  reg        [3:0]    _zz_PcPlugin_logic_harts_0_aggregator_oh_4;
  wire       [3:0]    PcPlugin_logic_harts_0_aggregator_oh;
  (* keep , syn_keep *) wire       [38:0]   PcPlugin_logic_harts_0_aggregator_target /* synthesis syn_keep = 1 */ ;
  wire                PcPlugin_logic_harts_0_aggregator_fault;
  wire                _zz_PcPlugin_logic_harts_0_aggregator_target;
  wire                _zz_PcPlugin_logic_harts_0_aggregator_target_1;
  wire                _zz_PcPlugin_logic_harts_0_aggregator_target_2;
  wire                _zz_PcPlugin_logic_harts_0_aggregator_fault_1;
  wire                when_PcPlugin_l80;
  wire                PcPlugin_logic_harts_0_holdComb;
  reg                 PcPlugin_logic_harts_0_holdReg;
  wire                PcPlugin_logic_harts_0_output_valid;
  wire                PcPlugin_logic_harts_0_output_ready;
  reg        [38:0]   PcPlugin_logic_harts_0_output_payload_pc;
  wire                PcPlugin_logic_harts_0_output_payload_fault;
  wire                PcPlugin_logic_harts_0_output_fire;
  wire                PcPlugin_logic_holdHalter_doIt;
  wire                fetch_logic_ctrls_0_haltRequest_PcPlugin_l133;
  reg        [1:0]    FetchL1Plugin_logic_translationStorage_logic_sl_0_write_mask;
  reg        [4:0]    FetchL1Plugin_logic_translationStorage_logic_sl_0_write_address;
  reg                 FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_valid;
  reg        [21:0]   FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_virtualAddress;
  reg        [19:0]   FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_physicalAddress;
  reg                 FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowRead;
  reg                 FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowWrite;
  reg                 FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowExecute;
  reg                 FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowUser;
  reg                 FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_willIncrement;
  wire                FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_willClear;
  reg        [0:0]    FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_valueNext;
  reg        [0:0]    FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_value;
  wire                FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_willOverflowIfInc;
  wire                FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_willOverflow;
  reg        [0:0]    FetchL1Plugin_logic_translationStorage_logic_sl_1_write_mask;
  reg        [4:0]    FetchL1Plugin_logic_translationStorage_logic_sl_1_write_address;
  reg                 FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_valid;
  reg        [12:0]   FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_virtualAddress;
  reg        [10:0]   FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_physicalAddress;
  reg                 FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowRead;
  reg                 FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowWrite;
  reg                 FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowExecute;
  reg                 FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowUser;
  reg                 FetchL1Plugin_logic_translationStorage_logic_sl_1_allocId_willIncrement;
  wire                FetchL1Plugin_logic_translationStorage_logic_sl_1_allocId_willClear;
  wire                FetchL1Plugin_logic_translationStorage_logic_sl_1_allocId_willOverflowIfInc;
  wire                FetchL1Plugin_logic_translationStorage_logic_sl_1_allocId_willOverflow;
  reg        [2:0]    LsuPlugin_logic_translationStorage_logic_sl_0_write_mask;
  reg        [4:0]    LsuPlugin_logic_translationStorage_logic_sl_0_write_address;
  reg                 LsuPlugin_logic_translationStorage_logic_sl_0_write_data_valid;
  reg        [21:0]   LsuPlugin_logic_translationStorage_logic_sl_0_write_data_virtualAddress;
  reg        [19:0]   LsuPlugin_logic_translationStorage_logic_sl_0_write_data_physicalAddress;
  reg                 LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowRead;
  reg                 LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowWrite;
  reg                 LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowExecute;
  reg                 LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowUser;
  reg                 LsuPlugin_logic_translationStorage_logic_sl_0_allocId_willIncrement;
  wire                LsuPlugin_logic_translationStorage_logic_sl_0_allocId_willClear;
  reg        [1:0]    LsuPlugin_logic_translationStorage_logic_sl_0_allocId_valueNext;
  reg        [1:0]    LsuPlugin_logic_translationStorage_logic_sl_0_allocId_value;
  wire                LsuPlugin_logic_translationStorage_logic_sl_0_allocId_willOverflowIfInc;
  wire                LsuPlugin_logic_translationStorage_logic_sl_0_allocId_willOverflow;
  reg        [0:0]    LsuPlugin_logic_translationStorage_logic_sl_1_write_mask;
  reg        [4:0]    LsuPlugin_logic_translationStorage_logic_sl_1_write_address;
  reg                 LsuPlugin_logic_translationStorage_logic_sl_1_write_data_valid;
  reg        [12:0]   LsuPlugin_logic_translationStorage_logic_sl_1_write_data_virtualAddress;
  reg        [10:0]   LsuPlugin_logic_translationStorage_logic_sl_1_write_data_physicalAddress;
  reg                 LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowRead;
  reg                 LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowWrite;
  reg                 LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowExecute;
  reg                 LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowUser;
  reg                 LsuPlugin_logic_translationStorage_logic_sl_1_allocId_willIncrement;
  wire                LsuPlugin_logic_translationStorage_logic_sl_1_allocId_willClear;
  wire                LsuPlugin_logic_translationStorage_logic_sl_1_allocId_willOverflowIfInc;
  wire                LsuPlugin_logic_translationStorage_logic_sl_1_allocId_willOverflow;
  wire                MmuPlugin_logic_isMachine;
  wire                MmuPlugin_logic_isSupervisor;
  wire                MmuPlugin_logic_isUser;
  wire                when_MmuPlugin_l277;
  wire                when_MmuPlugin_l279;
  wire       [4:0]    LsuPlugin_logic_onAddress0_translationPort_logic_read_0_readAddress;
  wire       [46:0]   _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_valid;
  wire       [46:0]   _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_valid;
  wire       [46:0]   _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_valid;
  wire       [4:0]    LsuPlugin_logic_onAddress0_translationPort_logic_read_1_readAddress;
  wire       [28:0]   _zz_execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_valid;
  wire       [3:0]    LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits;
  wire                LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hit;
  wire       [3:0]    _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_0;
  wire                LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_0;
  wire                LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_1;
  wire                LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_2;
  wire                LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_3;
  reg        [3:0]    _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_oh;
  wire                LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_range_0_to_1;
  wire                LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_range_0_to_2;
  wire       [3:0]    LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_oh;
  wire                _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute;
  wire                _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_1;
  wire                _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_2;
  wire                _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_3;
  wire                LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute;
  wire                LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowRead;
  wire                LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowWrite;
  wire                LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowUser;
  wire       [31:0]   LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated;
  reg                 LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_requireMmuLockup;
  wire       [4:0]    FetchL1Plugin_logic_translationPort_logic_read_0_readAddress;
  wire       [46:0]   _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_valid;
  wire       [46:0]   _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_valid;
  wire       [4:0]    FetchL1Plugin_logic_translationPort_logic_read_1_readAddress;
  wire       [28:0]   _zz_fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_valid;
  wire       [2:0]    FetchL1Plugin_logic_translationPort_logic_ctrl_hits;
  wire                FetchL1Plugin_logic_translationPort_logic_ctrl_hit;
  wire       [2:0]    _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_0;
  wire                FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_0;
  wire                FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_1;
  wire                FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_2;
  reg        [2:0]    _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_oh;
  wire                FetchL1Plugin_logic_translationPort_logic_ctrl_hits_range_0_to_1;
  wire       [2:0]    FetchL1Plugin_logic_translationPort_logic_ctrl_oh;
  wire                _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute;
  wire                _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_1;
  wire                _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_2;
  wire                FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute;
  wire                FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowRead;
  wire                FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowWrite;
  wire                FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowUser;
  wire       [31:0]   FetchL1Plugin_logic_translationPort_logic_ctrl_lineTranslated;
  reg                 FetchL1Plugin_logic_translationPort_logic_ctrl_requireMmuLockup;
  wire                MmuPlugin_logic_refill_wantExit;
  reg                 MmuPlugin_logic_refill_wantStart;
  wire                MmuPlugin_logic_refill_wantKill;
  wire                MmuPlugin_logic_refill_busy;
  reg        [38:0]   MmuPlugin_logic_refill_virtual;
  reg                 MmuPlugin_logic_refill_cacheRefillAny;
  reg                 MmuPlugin_logic_refill_cacheRefillAnySet;
  reg        [0:0]    MmuPlugin_logic_refill_portOhReg;
  reg        [1:0]    MmuPlugin_logic_refill_storageOhReg;
  reg                 MmuPlugin_logic_refill_storageEnable;
  wire                MmuPlugin_logic_refill_events_onStorage_0_waiting;
  wire                MmuPlugin_logic_refill_events_onStorage_1_waiting;
  reg        [31:0]   MmuPlugin_logic_refill_load_address;
  wire                MmuPlugin_logic_accessBus_rsp_toStream_valid;
  reg                 MmuPlugin_logic_accessBus_rsp_toStream_ready;
  wire       [63:0]   MmuPlugin_logic_accessBus_rsp_toStream_payload_data;
  wire                MmuPlugin_logic_accessBus_rsp_toStream_payload_error;
  wire                MmuPlugin_logic_accessBus_rsp_toStream_payload_redo;
  wire                MmuPlugin_logic_accessBus_rsp_toStream_payload_waitAny;
  wire                MmuPlugin_logic_refill_load_rsp_valid;
  reg                 MmuPlugin_logic_refill_load_rsp_ready;
  wire       [63:0]   MmuPlugin_logic_refill_load_rsp_payload_data;
  wire                MmuPlugin_logic_refill_load_rsp_payload_error;
  wire                MmuPlugin_logic_refill_load_rsp_payload_redo;
  wire                MmuPlugin_logic_refill_load_rsp_payload_waitAny;
  reg                 MmuPlugin_logic_accessBus_rsp_toStream_rValid;
  reg        [63:0]   MmuPlugin_logic_accessBus_rsp_toStream_rData_data;
  reg                 MmuPlugin_logic_accessBus_rsp_toStream_rData_error;
  reg                 MmuPlugin_logic_accessBus_rsp_toStream_rData_redo;
  reg                 MmuPlugin_logic_accessBus_rsp_toStream_rData_waitAny;
  wire                when_Stream_l477_2;
  wire       [63:0]   MmuPlugin_logic_refill_load_readed;
  wire                when_MmuPlugin_l400;
  wire                MmuPlugin_logic_refill_load_flags_V;
  wire                MmuPlugin_logic_refill_load_flags_R;
  wire                MmuPlugin_logic_refill_load_flags_W;
  wire                MmuPlugin_logic_refill_load_flags_X;
  wire                MmuPlugin_logic_refill_load_flags_U;
  wire                MmuPlugin_logic_refill_load_flags_G;
  wire                MmuPlugin_logic_refill_load_flags_A;
  wire                MmuPlugin_logic_refill_load_flags_D;
  wire       [63:0]   _zz_MmuPlugin_logic_refill_load_flags_V;
  wire                MmuPlugin_logic_refill_load_leaf;
  wire                MmuPlugin_logic_refill_load_reservedFault;
  reg                 MmuPlugin_logic_refill_load_exception;
  reg        [55:0]   MmuPlugin_logic_refill_load_levelToPhysicalAddress_0;
  reg        [55:0]   MmuPlugin_logic_refill_load_levelToPhysicalAddress_1;
  reg        [55:0]   MmuPlugin_logic_refill_load_levelToPhysicalAddress_2;
  wire                MmuPlugin_logic_refill_load_levelException_0;
  reg                 MmuPlugin_logic_refill_load_levelException_1;
  reg                 MmuPlugin_logic_refill_load_levelException_2;
  reg        [31:0]   MmuPlugin_logic_refill_load_nextLevelBase;
  wire                when_MmuPlugin_l421;
  wire                when_MmuPlugin_l421_1;
  wire                when_MmuPlugin_l421_2;
  wire                MmuPlugin_logic_refill_fetch_0_pteFault;
  wire                MmuPlugin_logic_refill_fetch_0_leafAccessFault;
  wire                MmuPlugin_logic_refill_fetch_0_pageFault;
  wire                MmuPlugin_logic_refill_fetch_0_accessFault;
  wire                MmuPlugin_logic_refill_fetch_1_pteFault;
  wire                MmuPlugin_logic_refill_fetch_1_leafAccessFault;
  wire                MmuPlugin_logic_refill_fetch_1_pageFault;
  wire                MmuPlugin_logic_refill_fetch_1_accessFault;
  wire                MmuPlugin_logic_refill_fetch_2_pteFault;
  wire                MmuPlugin_logic_refill_fetch_2_leafAccessFault;
  wire                MmuPlugin_logic_refill_fetch_2_pageFault;
  wire                MmuPlugin_logic_refill_fetch_2_accessFault;
  reg        [4:0]    MmuPlugin_logic_invalidate_counter;
  reg                 MmuPlugin_logic_invalidate_busy;
  wire                when_MmuPlugin_l565;
  wire                when_MmuPlugin_l579;
  reg        [11:0]   HistoryPlugin_logic_onFetch_value;
  reg        [11:0]   HistoryPlugin_logic_onFetch_valueNext;
  wire                HistoryPlugin_logic_onFetch_ports_0_valid;
  wire       [11:0]   HistoryPlugin_logic_onFetch_ports_0_payload_history;
  wire                HistoryPlugin_logic_onFetch_ports_1_valid;
  wire       [11:0]   HistoryPlugin_logic_onFetch_ports_1_payload_history;
  wire                HistoryPlugin_logic_onFetch_ports_2_valid;
  wire       [11:0]   HistoryPlugin_logic_onFetch_ports_2_payload_history;
  reg                 PerformanceCounterPlugin_logic_interrupt_ip;
  reg                 PerformanceCounterPlugin_logic_interrupt_ie;
  reg                 PerformanceCounterPlugin_logic_interrupt_sup_deleg;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_0;
  wire       [0:0]    PerformanceCounterPlugin_logic_events_sums_0;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_1;
  wire       [0:0]    PerformanceCounterPlugin_logic_events_sums_1;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_2;
  wire       [0:0]    PerformanceCounterPlugin_logic_events_sums_2;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_3;
  wire       [0:0]    PerformanceCounterPlugin_logic_events_sums_3;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_4;
  wire       [0:0]    PerformanceCounterPlugin_logic_events_sums_4;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_5;
  wire       [0:0]    PerformanceCounterPlugin_logic_events_sums_5;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_6;
  wire       [0:0]    PerformanceCounterPlugin_logic_events_sums_6;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_7;
  wire       [0:0]    PerformanceCounterPlugin_logic_events_sums_7;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_8;
  wire       [0:0]    PerformanceCounterPlugin_logic_events_sums_8;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_9;
  wire       [0:0]    PerformanceCounterPlugin_logic_events_sums_9;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_10;
  wire       [0:0]    PerformanceCounterPlugin_logic_events_sums_10;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_11;
  wire       [0:0]    PerformanceCounterPlugin_logic_events_sums_11;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_12;
  wire       [0:0]    PerformanceCounterPlugin_logic_events_sums_12;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_13;
  wire       [0:0]    PerformanceCounterPlugin_logic_events_sums_13;
  wire                PerformanceCounterPlugin_logic_fsm_wantExit;
  reg                 PerformanceCounterPlugin_logic_fsm_wantStart;
  wire                PerformanceCounterPlugin_logic_fsm_wantKill;
  wire                PerformanceCounterPlugin_logic_fsm_flusherCmd_valid;
  reg                 PerformanceCounterPlugin_logic_fsm_flusherCmd_ready;
  wire       [1:0]    PerformanceCounterPlugin_logic_fsm_flusherCmd_payload_oh;
  reg                 PerformanceCounterPlugin_logic_fsm_csrWriteCmd_valid;
  reg                 PerformanceCounterPlugin_logic_fsm_csrWriteCmd_ready;
  wire       [1:0]    PerformanceCounterPlugin_logic_fsm_csrWriteCmd_payload_address;
  wire                PerformanceCounterPlugin_logic_fsm_csrReadCmd_valid;
  reg                 PerformanceCounterPlugin_logic_fsm_csrReadCmd_ready;
  wire       [1:0]    PerformanceCounterPlugin_logic_fsm_csrReadCmd_payload_address;
  reg                 PerformanceCounterPlugin_logic_fsm_cmd_flusher;
  reg        [1:0]    PerformanceCounterPlugin_logic_fsm_cmd_oh;
  wire                _zz_PerformanceCounterPlugin_logic_fsm_cmd_address;
  wire                _zz_PerformanceCounterPlugin_logic_fsm_cmd_address_1;
  wire       [3:0]    PerformanceCounterPlugin_logic_fsm_cmd_address;
  wire                PerformanceCounterPlugin_logic_fsm_done;
  reg        [63:0]   PerformanceCounterPlugin_logic_fsm_ramReaded;
  reg                 PerformanceCounterPlugin_logic_fsm_carry;
  reg        [7:0]    PerformanceCounterPlugin_logic_fsm_counterReaded;
  wire       [63:0]   PerformanceCounterPlugin_logic_fsm_calc_a;
  wire       [7:0]    PerformanceCounterPlugin_logic_fsm_calc_b;
  wire       [64:0]   PerformanceCounterPlugin_logic_fsm_calc_sum;
  wire       [1:0]    PerformanceCounterPlugin_logic_fsm_idleCsrAddress;
  reg                 PerformanceCounterPlugin_logic_fsm_holdCsrWrite;
  wire       [1:0]    PerformanceCounterPlugin_logic_flusher_hits;
  wire                PerformanceCounterPlugin_logic_flusher_hit;
  wire       [1:0]    PerformanceCounterPlugin_logic_flusher_hits_ohFirst_input;
  wire       [1:0]    PerformanceCounterPlugin_logic_flusher_hits_ohFirst_masked;
  wire       [1:0]    PerformanceCounterPlugin_logic_flusher_oh;
  wire       [1:0]    PerformanceCounterPlugin_logic_csrDecode_addr;
  reg                 PerformanceCounterPlugin_logic_csrDecode_mok;
  reg                 PerformanceCounterPlugin_logic_csrDecode_sok;
  wire                PerformanceCounterPlugin_logic_csrDecode_privOk;
  reg                 PerformanceCounterPlugin_logic_csrRead_fired;
  wire                PerformanceCounterPlugin_logic_fsm_csrReadCmd_fire;
  wire                PerformanceCounterPlugin_logic_csrRead_requested;
  wire                when_PerformanceCounterPlugin_l342;
  reg                 PerformanceCounterPlugin_logic_csrWrite_fired;
  wire                PerformanceCounterPlugin_logic_fsm_csrWriteCmd_fire;
  wire                fetch_logic_flushes_0_doIt;
  wire                fetch_logic_ctrls_1_throwWhen_FetchPipelinePlugin_l48;
  wire                fetch_logic_flushes_1_doIt;
  wire                fetch_logic_ctrls_2_forgetsSingleRequest_FetchPipelinePlugin_l50;
  wire                CsrAccessPlugin_logic_fsm_wantExit;
  reg                 CsrAccessPlugin_logic_fsm_wantStart;
  wire                CsrAccessPlugin_logic_fsm_wantKill;
  reg                 REG_CSR_768;
  reg                 REG_CSR_256;
  reg                 REG_CSR_384;
  reg                 REG_CSR_944;
  reg                 REG_CSR_928;
  reg                 REG_CSR_945;
  reg                 REG_CSR_946;
  reg                 REG_CSR_947;
  reg                 REG_CSR_PmpPlugin_logic_allFilter;
  reg                 REG_CSR_794;
  reg                 REG_CSR_1952;
  reg                 REG_CSR_1953;
  reg                 REG_CSR_1954;
  reg                 REG_CSR_3857;
  reg                 REG_CSR_3858;
  reg                 REG_CSR_3859;
  reg                 REG_CSR_3860;
  reg                 REG_CSR_769;
  reg                 REG_CSR_834;
  reg                 REG_CSR_836;
  reg                 REG_CSR_772;
  reg                 REG_CSR_770;
  reg                 REG_CSR_771;
  reg                 REG_CSR_4016;
  reg                 REG_CSR_774;
  reg                 REG_CSR_322;
  reg                 REG_CSR_778;
  reg                 REG_CSR_260;
  reg                 REG_CSR_324;
  reg                 REG_CSR_3504;
  reg                 REG_CSR_3073;
  reg                 REG_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_tvecFilter;
  reg                 REG_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_epcFilter;
  reg                 REG_CSR_262;
  reg                 REG_CSR_800;
  reg                 REG_CSR_UNAMED_0;
  reg                 REG_CSR_266;
  reg                 REG_CSR_CsrRamPlugin_csrMapper_selFilter;
  reg                 REG_CSR_PerformanceCounterPlugin_logic_csrFilter;
  reg                 REG_CSR_CsrAccessPlugin_logic_trapNextOnWriteFilter;
  reg                 CsrAccessPlugin_logic_fsm_interface_read;
  reg                 CsrAccessPlugin_logic_fsm_interface_write;
  wire       [63:0]   CsrAccessPlugin_logic_fsm_interface_rs1;
  reg        [63:0]   CsrAccessPlugin_logic_fsm_interface_aluInput;
  reg        [63:0]   CsrAccessPlugin_logic_fsm_interface_csrValue;
  reg        [63:0]   CsrAccessPlugin_logic_fsm_interface_onWriteBits;
  wire       [15:0]   CsrAccessPlugin_logic_fsm_interface_uopId;
  wire       [31:0]   CsrAccessPlugin_logic_fsm_interface_uop;
  wire                CsrAccessPlugin_logic_fsm_interface_doImm;
  wire                CsrAccessPlugin_logic_fsm_interface_doMask;
  wire                CsrAccessPlugin_logic_fsm_interface_doClear;
  wire       [4:0]    CsrAccessPlugin_logic_fsm_interface_rdPhys;
  wire                CsrAccessPlugin_logic_fsm_interface_rdEnable;
  reg                 CsrAccessPlugin_logic_fsm_interface_fire;
  wire       [11:0]   CsrAccessPlugin_logic_fsm_inject_csrAddress;
  wire                CsrAccessPlugin_logic_fsm_inject_immZero;
  wire                CsrAccessPlugin_logic_fsm_inject_srcZero;
  wire                CsrAccessPlugin_logic_fsm_inject_csrWrite;
  wire                CsrAccessPlugin_logic_fsm_inject_csrRead;
  wire                COMB_CSR_768;
  wire                COMB_CSR_256;
  wire                COMB_CSR_384;
  wire                COMB_CSR_944;
  wire                COMB_CSR_928;
  wire                COMB_CSR_945;
  wire                COMB_CSR_946;
  wire                COMB_CSR_947;
  wire                COMB_CSR_PmpPlugin_logic_allFilter;
  wire                COMB_CSR_794;
  wire                COMB_CSR_1952;
  wire                COMB_CSR_1953;
  wire                COMB_CSR_1954;
  wire                COMB_CSR_3857;
  wire                COMB_CSR_3858;
  wire                COMB_CSR_3859;
  wire                COMB_CSR_3860;
  wire                COMB_CSR_769;
  wire                COMB_CSR_834;
  wire                COMB_CSR_836;
  wire                COMB_CSR_772;
  wire                COMB_CSR_770;
  wire                COMB_CSR_771;
  wire                COMB_CSR_4016;
  wire                COMB_CSR_774;
  wire                COMB_CSR_322;
  wire                COMB_CSR_778;
  wire                COMB_CSR_260;
  wire                COMB_CSR_324;
  wire                COMB_CSR_3504;
  wire                COMB_CSR_3073;
  wire                COMB_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_tvecFilter;
  wire                COMB_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_epcFilter;
  wire                COMB_CSR_262;
  wire                COMB_CSR_800;
  wire                COMB_CSR_UNAMED_1;
  wire                COMB_CSR_266;
  wire                COMB_CSR_CsrRamPlugin_csrMapper_selFilter;
  wire                COMB_CSR_PerformanceCounterPlugin_logic_csrFilter;
  wire                COMB_CSR_CsrAccessPlugin_logic_trapNextOnWriteFilter;
  wire                CsrAccessPlugin_logic_fsm_inject_implemented;
  wire                CsrAccessPlugin_logic_fsm_inject_onDecodeDo;
  wire                when_CsrAccessPlugin_l157;
  wire                when_MmuPlugin_l223;
  wire                when_CsrAccessPlugin_l157_1;
  wire                when_CsrAccessPlugin_l157_2;
  wire                when_CsrService_l121;
  wire                when_CsrAccessPlugin_l157_3;
  wire                when_CsrService_l121_1;
  wire                when_CsrAccessPlugin_l157_4;
  wire                when_CsrService_l121_2;
  wire                when_CsrAccessPlugin_l157_5;
  wire                when_CsrService_l121_3;
  wire                when_CsrAccessPlugin_l157_6;
  wire                when_CsrService_l198;
  wire                when_CsrService_l199;
  wire                when_CsrAccessPlugin_l157_7;
  wire                when_CsrService_l121_4;
  wire                when_CsrAccessPlugin_l157_8;
  wire                when_CsrService_l121_5;
  wire                when_CsrAccessPlugin_l157_9;
  wire                when_PerformanceCounterPlugin_l327;
  wire                when_PerformanceCounterPlugin_l328;
  wire                when_CsrAccessPlugin_l157_10;
  wire                CsrAccessPlugin_logic_fsm_inject_trap;
  reg                 CsrAccessPlugin_logic_fsm_inject_unfreeze;
  wire                CsrAccessPlugin_logic_fsm_inject_freeze;
  reg                 CsrAccessPlugin_logic_fsm_inject_flushReg;
  wire                when_CsrAccessPlugin_l199;
  reg                 CsrAccessPlugin_logic_fsm_inject_sampled;
  reg                 CsrAccessPlugin_logic_fsm_inject_trapReg;
  reg                 CsrAccessPlugin_logic_fsm_inject_busTrapReg;
  reg        [3:0]    CsrAccessPlugin_logic_fsm_inject_busTrapCodeReg;
  reg                 CsrAccessPlugin_logic_fsm_readLogic_onReadsDo;
  reg                 CsrAccessPlugin_logic_fsm_readLogic_onReadsFireDo;
  wire                when_CsrAccessPlugin_l258;
  wire       [63:0]   CsrAccessPlugin_logic_fsm_readLogic_csrValue;
  wire                when_CsrAccessPlugin_l285;
  wire       [63:0]   CsrAccessPlugin_logic_fsm_writeLogic_alu_mask;
  wire       [63:0]   CsrAccessPlugin_logic_fsm_writeLogic_alu_masked;
  wire       [63:0]   CsrAccessPlugin_logic_fsm_writeLogic_alu_result;
  reg                 CsrAccessPlugin_logic_fsm_writeLogic_onWritesDo;
  reg                 CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo;
  wire                when_CsrAccessPlugin_l352;
  wire       [1:0]    switch_PrivilegedPlugin_l581;
  wire                when_CsrAccessPlugin_l352_1;
  wire                when_CsrAccessPlugin_l359;
  wire                when_CsrAccessPlugin_l352_2;
  wire                when_CsrAccessPlugin_l359_1;
  wire                when_CsrAccessPlugin_l352_3;
  wire                when_CsrAccessPlugin_l352_4;
  wire                when_CsrAccessPlugin_l359_2;
  wire                when_CsrAccessPlugin_l352_5;
  wire                when_CsrAccessPlugin_l359_3;
  wire                when_CsrAccessPlugin_l352_6;
  wire                when_CsrAccessPlugin_l359_4;
  wire                when_CsrAccessPlugin_l352_7;
  wire                when_CsrAccessPlugin_l352_8;
  wire                when_CsrAccessPlugin_l352_9;
  wire                when_CsrAccessPlugin_l352_10;
  wire                when_CsrAccessPlugin_l352_11;
  wire                when_CsrAccessPlugin_l352_12;
  wire                when_CsrAccessPlugin_l352_13;
  wire                when_CsrAccessPlugin_l352_14;
  wire                when_CsrAccessPlugin_l352_15;
  wire                when_CsrAccessPlugin_l352_16;
  wire                when_CsrAccessPlugin_l352_17;
  wire                when_CsrAccessPlugin_l349;
  wire                when_CsrAccessPlugin_l349_1;
  wire                when_CsrAccessPlugin_l352_18;
  wire                when_CsrAccessPlugin_l352_19;
  wire                when_CsrAccessPlugin_l352_20;
  wire                when_CsrAccessPlugin_l349_2;
  wire                when_CsrAccessPlugin_l349_3;
  wire                when_PerformanceCounterPlugin_l357;
  wire                when_PerformanceCounterPlugin_l359;
  wire       [3:0]    CsrRamPlugin_logic_writeLogic_hits;
  wire                CsrRamPlugin_logic_writeLogic_hit;
  wire       [3:0]    CsrRamPlugin_logic_writeLogic_hits_ohFirst_input;
  wire       [3:0]    CsrRamPlugin_logic_writeLogic_hits_ohFirst_masked;
  wire       [3:0]    CsrRamPlugin_logic_writeLogic_oh;
  wire                CsrRamPlugin_logic_writeLogic_port_valid;
  wire       [3:0]    CsrRamPlugin_logic_writeLogic_port_payload_address;
  wire       [63:0]   CsrRamPlugin_logic_writeLogic_port_payload_data;
  wire                _zz_PerformanceCounterPlugin_logic_writePort_ready;
  wire                _zz_TrapPlugin_logic_harts_0_crsPorts_write_ready;
  wire                _zz_CsrRamPlugin_csrMapper_write_ready;
  wire                _zz_CsrRamPlugin_setup_initPort_ready;
  wire       [2:0]    CsrRamPlugin_logic_readLogic_hits;
  wire                CsrRamPlugin_logic_readLogic_hit;
  wire       [2:0]    CsrRamPlugin_logic_readLogic_hits_ohFirst_input;
  wire       [2:0]    CsrRamPlugin_logic_readLogic_hits_ohFirst_masked;
  wire       [2:0]    CsrRamPlugin_logic_readLogic_oh;
  wire                _zz_CsrRamPlugin_logic_readLogic_sel;
  wire                _zz_CsrRamPlugin_logic_readLogic_sel_1;
  wire       [1:0]    CsrRamPlugin_logic_readLogic_sel;
  wire                CsrRamPlugin_logic_readLogic_port_cmd_valid;
  wire       [3:0]    CsrRamPlugin_logic_readLogic_port_cmd_payload;
  wire       [63:0]   CsrRamPlugin_logic_readLogic_port_rsp;
  reg        [2:0]    CsrRamPlugin_logic_readLogic_ohReg;
  reg                 CsrRamPlugin_logic_readLogic_busy;
  reg        [4:0]    CsrRamPlugin_logic_flush_counter;
  wire                CsrRamPlugin_logic_flush_done;
  wire                execute_lane0_bypasser_integer_RS1_port_valid;
  wire       [4:0]    execute_lane0_bypasser_integer_RS1_port_address;
  wire       [63:0]   execute_lane0_bypasser_integer_RS1_port_data;
  reg        [4:0]    execute_lane0_bypasser_integer_RS1_bypassEnables;
  wire       [4:0]    _zz_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0;
  wire                execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0;
  wire                execute_lane0_bypasser_integer_RS1_bypassEnables_bools_1;
  wire                execute_lane0_bypasser_integer_RS1_bypassEnables_bools_2;
  wire                execute_lane0_bypasser_integer_RS1_bypassEnables_bools_3;
  wire                execute_lane0_bypasser_integer_RS1_bypassEnables_bools_4;
  reg        [4:0]    _zz_execute_lane0_bypasser_integer_RS1_sel;
  wire                execute_lane0_bypasser_integer_RS1_bypassEnables_range_0_to_1;
  wire                execute_lane0_bypasser_integer_RS1_bypassEnables_range_0_to_2;
  wire                execute_lane0_bypasser_integer_RS1_bypassEnables_range_0_to_3;
  wire       [4:0]    execute_lane0_bypasser_integer_RS1_sel;
  wire       [3:0]    _zz_execute_ctrl1_down_integer_RS1_lane0;
  (* keep , syn_keep *) reg        [63:0]   _zz_execute_ctrl1_down_integer_RS1_lane0_1 /* synthesis syn_keep = 1 */ ;
  wire                when_ExecuteLanePlugin_l196;
  wire                execute_lane0_bypasser_integer_RS2_port_valid;
  wire       [4:0]    execute_lane0_bypasser_integer_RS2_port_address;
  wire       [63:0]   execute_lane0_bypasser_integer_RS2_port_data;
  reg        [4:0]    execute_lane0_bypasser_integer_RS2_bypassEnables;
  wire       [4:0]    _zz_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0;
  wire                execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0;
  wire                execute_lane0_bypasser_integer_RS2_bypassEnables_bools_1;
  wire                execute_lane0_bypasser_integer_RS2_bypassEnables_bools_2;
  wire                execute_lane0_bypasser_integer_RS2_bypassEnables_bools_3;
  wire                execute_lane0_bypasser_integer_RS2_bypassEnables_bools_4;
  reg        [4:0]    _zz_execute_lane0_bypasser_integer_RS2_sel;
  wire                execute_lane0_bypasser_integer_RS2_bypassEnables_range_0_to_1;
  wire                execute_lane0_bypasser_integer_RS2_bypassEnables_range_0_to_2;
  wire                execute_lane0_bypasser_integer_RS2_bypassEnables_range_0_to_3;
  wire       [4:0]    execute_lane0_bypasser_integer_RS2_sel;
  wire       [3:0]    _zz_execute_ctrl1_down_integer_RS2_lane0;
  (* keep , syn_keep *) reg        [63:0]   _zz_execute_ctrl1_down_integer_RS2_lane0_1 /* synthesis syn_keep = 1 */ ;
  wire                when_ExecuteLanePlugin_l196_1;
  wire                execute_lane0_logic_completions_onCtrl_0_port_valid;
  wire       [15:0]   execute_lane0_logic_completions_onCtrl_0_port_payload_uopId;
  wire                execute_lane0_logic_completions_onCtrl_0_port_payload_trap;
  wire                execute_lane0_logic_completions_onCtrl_0_port_payload_commit;
  wire                execute_lane0_logic_completions_onCtrl_1_port_valid;
  wire       [15:0]   execute_lane0_logic_completions_onCtrl_1_port_payload_uopId;
  wire                execute_lane0_logic_completions_onCtrl_1_port_payload_trap;
  wire                execute_lane0_logic_completions_onCtrl_1_port_payload_commit;
  wire                execute_lane0_logic_completions_onCtrl_2_port_valid;
  wire       [15:0]   execute_lane0_logic_completions_onCtrl_2_port_payload_uopId;
  wire                execute_lane0_logic_completions_onCtrl_2_port_payload_trap;
  wire                execute_lane0_logic_completions_onCtrl_2_port_payload_commit;
  wire       [31:0]   execute_lane0_logic_decoding_decodingBits;
  wire                _zz_execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0_1;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0_2;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_1;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_2;
  wire                _zz_execute_ctrl1_down_AguPlugin_LOAD_lane0;
  wire                _zz_execute_ctrl1_down_BYPASSED_AT_3_lane0;
  wire                _zz_execute_ctrl1_down_AguPlugin_ATOMIC_lane0;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_1;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_2;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_3;
  wire                _zz_execute_ctrl1_down_BYPASSED_AT_3_lane0_1;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_3;
  wire                _zz_execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0;
  wire                _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0;
  wire                _zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0;
  wire                _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0;
  wire       [1:0]    _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  wire       [1:0]    _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1;
  wire       [1:0]    _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2;
  wire                _zz_execute_ctrl1_down_BYPASSED_AT_3_lane0_2;
  wire                _zz_execute_ctrl1_down_RsUnsignedPlugin_IS_W_lane0;
  wire                _zz_execute_ctrl1_down_AguPlugin_STORE_lane0;
  wire       [1:0]    _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0;
  wire       [1:0]    _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_1;
  wire       [1:0]    _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_2;
  wire                _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0;
  wire                _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0;
  wire       [2:0]    _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1;
  wire       [2:0]    _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2;
  wire       [2:0]    _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_3;
  wire                when_ExecuteLanePlugin_l306;
  wire                when_ExecuteLanePlugin_l306_1;
  wire                when_ExecuteLanePlugin_l306_2;
  wire                when_ExecuteLanePlugin_l306_3;
  wire                when_ExecuteLanePlugin_l306_4;
  wire                WhiteboxerPlugin_logic_csr_port_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_csr_port_payload_uopId;
  wire       [11:0]   WhiteboxerPlugin_logic_csr_port_payload_address;
  wire       [63:0]   WhiteboxerPlugin_logic_csr_port_payload_write;
  wire       [63:0]   WhiteboxerPlugin_logic_csr_port_payload_read;
  wire                WhiteboxerPlugin_logic_csr_port_payload_writeDone;
  wire                WhiteboxerPlugin_logic_csr_port_payload_readDone;
  wire                WhiteboxerPlugin_logic_rfWrites_ports_0_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_rfWrites_ports_0_payload_uopId;
  wire       [63:0]   WhiteboxerPlugin_logic_rfWrites_ports_0_payload_data;
  wire                WhiteboxerPlugin_logic_rfWrites_ports_1_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_rfWrites_ports_1_payload_uopId;
  wire       [63:0]   WhiteboxerPlugin_logic_rfWrites_ports_1_payload_data;
  wire                WhiteboxerPlugin_logic_rfWrites_ports_2_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_rfWrites_ports_2_payload_uopId;
  wire       [63:0]   WhiteboxerPlugin_logic_rfWrites_ports_2_payload_data;
  wire                WhiteboxerPlugin_logic_completions_ports_0_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_completions_ports_0_payload_uopId;
  wire                WhiteboxerPlugin_logic_completions_ports_0_payload_trap;
  wire                WhiteboxerPlugin_logic_completions_ports_0_payload_commit;
  wire                WhiteboxerPlugin_logic_completions_ports_1_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_completions_ports_1_payload_uopId;
  wire                WhiteboxerPlugin_logic_completions_ports_1_payload_trap;
  wire                WhiteboxerPlugin_logic_completions_ports_1_payload_commit;
  wire                WhiteboxerPlugin_logic_completions_ports_2_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_completions_ports_2_payload_uopId;
  wire                WhiteboxerPlugin_logic_completions_ports_2_payload_trap;
  wire                WhiteboxerPlugin_logic_completions_ports_2_payload_commit;
  wire                WhiteboxerPlugin_logic_completions_ports_3_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_completions_ports_3_payload_uopId;
  wire                WhiteboxerPlugin_logic_completions_ports_3_payload_trap;
  wire                WhiteboxerPlugin_logic_completions_ports_3_payload_commit;
  wire                WhiteboxerPlugin_logic_commits_ports_0_oh_0;
  wire                WhiteboxerPlugin_logic_commits_ports_0_valid;
  wire       [38:0]   WhiteboxerPlugin_logic_commits_ports_0_pc;
  wire       [31:0]   WhiteboxerPlugin_logic_commits_ports_0_uop;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_0_valid;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_0_payload_self;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_1_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_reschedules_flushes_1_payload_uopId;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_1_payload_self;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_2_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_reschedules_flushes_2_payload_uopId;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_2_payload_self;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_3_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_reschedules_flushes_3_payload_uopId;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_3_payload_self;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_4_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_reschedules_flushes_4_payload_uopId;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_4_payload_self;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_5_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_reschedules_flushes_5_payload_uopId;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_5_payload_self;
  wire                early0_BranchPlugin_logic_jumpLogic_learn_asFlow_valid;
  wire       [38:0]   early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_pcOnLastSlice;
  wire       [38:0]   early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_pcTarget;
  wire                early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_taken;
  wire                early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_isBranch;
  wire                early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_isPush;
  wire                early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_isPop;
  wire                early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_wasWrong;
  wire                early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_badPredictedTarget;
  wire       [11:0]   early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_history;
  wire       [15:0]   early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_uopId;
  wire       [1:0]    early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  wire                WhiteboxerPlugin_logic_prediction_learns_0_valid;
  wire       [38:0]   WhiteboxerPlugin_logic_prediction_learns_0_payload_pcOnLastSlice;
  wire       [38:0]   WhiteboxerPlugin_logic_prediction_learns_0_payload_pcTarget;
  wire                WhiteboxerPlugin_logic_prediction_learns_0_payload_taken;
  wire                WhiteboxerPlugin_logic_prediction_learns_0_payload_isBranch;
  wire                WhiteboxerPlugin_logic_prediction_learns_0_payload_isPush;
  wire                WhiteboxerPlugin_logic_prediction_learns_0_payload_isPop;
  wire                WhiteboxerPlugin_logic_prediction_learns_0_payload_wasWrong;
  wire                WhiteboxerPlugin_logic_prediction_learns_0_payload_badPredictedTarget;
  wire       [11:0]   WhiteboxerPlugin_logic_prediction_learns_0_payload_history;
  wire       [15:0]   WhiteboxerPlugin_logic_prediction_learns_0_payload_uopId;
  wire       [1:0]    WhiteboxerPlugin_logic_prediction_learns_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    WhiteboxerPlugin_logic_prediction_learns_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  wire                WhiteboxerPlugin_logic_loadExecute_fire;
  wire       [15:0]   WhiteboxerPlugin_logic_loadExecute_uopId;
  wire       [1:0]    WhiteboxerPlugin_logic_loadExecute_size;
  wire       [31:0]   WhiteboxerPlugin_logic_loadExecute_address;
  wire       [63:0]   WhiteboxerPlugin_logic_loadExecute_data;
  wire                WhiteboxerPlugin_logic_storeCommit_fire;
  wire       [15:0]   WhiteboxerPlugin_logic_storeCommit_uopId;
  wire       [11:0]   WhiteboxerPlugin_logic_storeCommit_storeId;
  wire       [1:0]    WhiteboxerPlugin_logic_storeCommit_size;
  wire       [31:0]   WhiteboxerPlugin_logic_storeCommit_address;
  wire       [63:0]   WhiteboxerPlugin_logic_storeCommit_data;
  wire                WhiteboxerPlugin_logic_storeCommit_amo;
  wire                WhiteboxerPlugin_logic_storeConditional_fire;
  wire       [15:0]   WhiteboxerPlugin_logic_storeConditional_uopId;
  wire                WhiteboxerPlugin_logic_storeConditional_miss;
  wire                WhiteboxerPlugin_logic_storeBroadcast_fire;
  wire       [11:0]   WhiteboxerPlugin_logic_storeBroadcast_storeId;
  wire                integer_RegFilePlugin_logic_writeMerges_0_bus_valid;
  wire       [4:0]    integer_RegFilePlugin_logic_writeMerges_0_bus_address;
  wire       [63:0]   integer_RegFilePlugin_logic_writeMerges_0_bus_data;
  wire       [15:0]   integer_RegFilePlugin_logic_writeMerges_0_bus_uopId;
  reg        [5:0]    integer_RegFilePlugin_logic_initalizer_counter;
  wire                integer_RegFilePlugin_logic_initalizer_done;
  wire                when_RegFilePlugin_l132;
  wire                integer_write_0_valid /* verilator public */ ;
  wire       [4:0]    integer_write_0_address /* verilator public */ ;
  wire       [63:0]   integer_write_0_data /* verilator public */ ;
  wire       [15:0]   integer_write_0_uopId /* verilator public */ ;
  wire       [0:0]    WhiteboxerPlugin_logic_wfi;
  wire                WhiteboxerPlugin_logic_perf_executeFreezed;
  wire                WhiteboxerPlugin_logic_perf_dispatchHazards;
  wire       [0:0]    WhiteboxerPlugin_logic_perf_candidatesCount;
  wire       [0:0]    WhiteboxerPlugin_logic_perf_dispatchFeedCount;
  reg                 _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_1;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_2;
  wire       [59:0]   WhiteboxerPlugin_logic_perf_executeFreezedCounter;
  reg                 _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_1;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_2;
  wire       [59:0]   WhiteboxerPlugin_logic_perf_dispatchHazardsCounter;
  wire                when_Utils_l598;
  reg                 _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_1;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_2;
  wire       [59:0]   WhiteboxerPlugin_logic_perf_candidatesCountCounters_0;
  wire                when_Utils_l598_1;
  reg                 _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_1;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_2;
  wire       [59:0]   WhiteboxerPlugin_logic_perf_candidatesCountCounters_1;
  wire                when_Utils_l598_2;
  reg                 _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_1;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_2;
  wire       [59:0]   WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0;
  wire                when_Utils_l598_3;
  reg                 _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_1;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_2;
  wire       [59:0]   WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1;
  wire                WhiteboxerPlugin_logic_trap_ports_0_valid;
  wire                WhiteboxerPlugin_logic_trap_ports_0_interrupt;
  wire       [3:0]    WhiteboxerPlugin_logic_trap_ports_0_cause;
  wire                fetch_logic_ctrls_2_up_forgetOne;
  wire                fetch_logic_ctrls_1_up_forgetOne;
  wire                when_CtrlLink_l191;
  wire                when_CtrlLink_l198;
  wire                when_StageLink_l71;
  wire                when_DecodePipelinePlugin_l70;
  reg        [1:0]    LsuPlugin_logic_flusher_stateReg;
  reg        [1:0]    LsuPlugin_logic_flusher_stateNext;
  wire                when_LsuPlugin_l368;
  wire                when_LsuPlugin_l376;
  wire                LsuPlugin_logic_flusher_onExit_IDLE;
  wire                LsuPlugin_logic_flusher_onExit_CMD;
  wire                LsuPlugin_logic_flusher_onExit_COMPLETION;
  wire                LsuPlugin_logic_flusher_onEntry_IDLE;
  wire                LsuPlugin_logic_flusher_onEntry_CMD;
  wire                LsuPlugin_logic_flusher_onEntry_COMPLETION;
  reg        [3:0]    TrapPlugin_logic_harts_0_trap_fsm_stateReg;
  reg        [3:0]    TrapPlugin_logic_harts_0_trap_fsm_stateNext;
  wire                when_TrapPlugin_l453;
  wire                when_TrapPlugin_l481;
  reg        [3:0]    _zz_TrapPlugin_logic_harts_0_crsPorts_write_address;
  reg        [3:0]    _zz_TrapPlugin_logic_harts_0_crsPorts_write_address_1;
  reg        [3:0]    _zz_TrapPlugin_logic_harts_0_crsPorts_read_address;
  wire                when_TrapPlugin_l615;
  reg        [3:0]    _zz_TrapPlugin_logic_harts_0_crsPorts_read_address_1;
  wire                when_TrapPlugin_l712;
  wire       [1:0]    switch_TrapPlugin_l713;
  wire                when_TrapPlugin_l555;
  wire       [2:0]    switch_TrapPlugin_l557;
  wire                when_TrapPlugin_l406;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onExit_RESET;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onExit_RUNNING;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onExit_COMPUTE;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onExit_TRAP_EPC;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onExit_TRAP_TVAL;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onExit_TRAP_TVEC;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onExit_TRAP_WAIT;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onExit_TRAP_APPLY;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onExit_XRET_EPC;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onExit_XRET_APPLY;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onExit_ATS_RSP;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onExit_JUMP;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onExit_LSU_FLUSH;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onExit_FETCH_FLUSH;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onEntry_RESET;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onEntry_RUNNING;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onEntry_COMPUTE;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onEntry_TRAP_EPC;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onEntry_TRAP_TVAL;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onEntry_TRAP_TVEC;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onEntry_TRAP_WAIT;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onEntry_TRAP_APPLY;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onEntry_XRET_EPC;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onEntry_XRET_APPLY;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onEntry_ATS_RSP;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onEntry_JUMP;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onEntry_LSU_FLUSH;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onEntry_FETCH_FLUSH;
  reg        [3:0]    MmuPlugin_logic_refill_stateReg;
  reg        [3:0]    MmuPlugin_logic_refill_stateNext;
  wire                when_MmuPlugin_l516;
  wire                when_MmuPlugin_l516_1;
  wire                when_MmuPlugin_l516_2;
  wire                when_MmuPlugin_l525;
  wire                when_MmuPlugin_l534;
  wire                when_MmuPlugin_l534_1;
  wire                _zz_55;
  wire                when_MmuPlugin_l505;
  wire                when_MmuPlugin_l505_1;
  wire                when_MmuPlugin_l505_2;
  wire                when_MmuPlugin_l505_3;
  wire                when_MmuPlugin_l505_4;
  wire                when_MmuPlugin_l505_5;
  wire                MmuPlugin_logic_refill_onExit_BOOT;
  wire                MmuPlugin_logic_refill_onExit_IDLE;
  wire                MmuPlugin_logic_refill_onExit_CMD_0;
  wire                MmuPlugin_logic_refill_onExit_CMD_1;
  wire                MmuPlugin_logic_refill_onExit_CMD_2;
  wire                MmuPlugin_logic_refill_onExit_RSP_0;
  wire                MmuPlugin_logic_refill_onExit_RSP_1;
  wire                MmuPlugin_logic_refill_onExit_RSP_2;
  wire                MmuPlugin_logic_refill_onExit_DONE_0;
  wire                MmuPlugin_logic_refill_onExit_DONE_1;
  wire                MmuPlugin_logic_refill_onExit_DONE_2;
  wire                MmuPlugin_logic_refill_onEntry_BOOT;
  wire                MmuPlugin_logic_refill_onEntry_IDLE;
  wire                MmuPlugin_logic_refill_onEntry_CMD_0;
  wire                MmuPlugin_logic_refill_onEntry_CMD_1;
  wire                MmuPlugin_logic_refill_onEntry_CMD_2;
  wire                MmuPlugin_logic_refill_onEntry_RSP_0;
  wire                MmuPlugin_logic_refill_onEntry_RSP_1;
  wire                MmuPlugin_logic_refill_onEntry_RSP_2;
  wire                MmuPlugin_logic_refill_onEntry_DONE_0;
  wire                MmuPlugin_logic_refill_onEntry_DONE_1;
  wire                MmuPlugin_logic_refill_onEntry_DONE_2;
  reg        [2:0]    PerformanceCounterPlugin_logic_fsm_stateReg;
  reg        [2:0]    PerformanceCounterPlugin_logic_fsm_stateNext;
  wire                when_PerformanceCounterPlugin_l271;
  wire                when_PerformanceCounterPlugin_l249;
  wire                when_PerformanceCounterPlugin_l255;
  wire                PerformanceCounterPlugin_logic_fsm_onExit_BOOT;
  wire                PerformanceCounterPlugin_logic_fsm_onExit_IDLE;
  wire                PerformanceCounterPlugin_logic_fsm_onExit_READ_LOW;
  wire                PerformanceCounterPlugin_logic_fsm_onExit_CALC_LOW;
  wire                PerformanceCounterPlugin_logic_fsm_onExit_CSR_WRITE;
  wire                PerformanceCounterPlugin_logic_fsm_onEntry_BOOT;
  wire                PerformanceCounterPlugin_logic_fsm_onEntry_IDLE;
  wire                PerformanceCounterPlugin_logic_fsm_onEntry_READ_LOW;
  wire                PerformanceCounterPlugin_logic_fsm_onEntry_CALC_LOW;
  wire                PerformanceCounterPlugin_logic_fsm_onEntry_CSR_WRITE;
  reg        [1:0]    CsrAccessPlugin_logic_fsm_stateReg;
  reg        [1:0]    CsrAccessPlugin_logic_fsm_stateNext;
  wire                when_CsrAccessPlugin_l302;
  wire                when_CsrAccessPlugin_l331;
  wire                when_CsrAccessPlugin_l214;
  wire                when_CsrAccessPlugin_l215;
  wire                when_CsrAccessPlugin_l227;
  wire                CsrAccessPlugin_logic_fsm_onExit_IDLE;
  wire                CsrAccessPlugin_logic_fsm_onExit_READ;
  wire                CsrAccessPlugin_logic_fsm_onExit_WRITE;
  wire                CsrAccessPlugin_logic_fsm_onExit_COMPLETION;
  wire                CsrAccessPlugin_logic_fsm_onEntry_IDLE;
  wire                CsrAccessPlugin_logic_fsm_onEntry_READ;
  wire                CsrAccessPlugin_logic_fsm_onEntry_WRITE;
  wire                CsrAccessPlugin_logic_fsm_onEntry_COMPLETION;
  `ifndef SYNTHESIS
  reg [79:0] execute_ctrl2_up_early0_EnvPlugin_OP_lane0_string;
  reg [31:0] execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane0_string;
  reg [39:0] execute_ctrl2_up_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string;
  reg [79:0] execute_ctrl1_down_early0_EnvPlugin_OP_lane0_string;
  reg [31:0] execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_string;
  reg [39:0] execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string;
  reg [31:0] execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0_string;
  reg [79:0] execute_ctrl2_down_early0_EnvPlugin_OP_lane0_string;
  reg [39:0] execute_ctrl2_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string;
  reg [95:0] LsuPlugin_logic_onAddress0_ls_port_payload_op_string;
  reg [95:0] LsuPlugin_logic_onAddress0_access_port_payload_op_string;
  reg [95:0] LsuPlugin_logic_onAddress0_flush_port_payload_op_string;
  reg [39:0] _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string;
  reg [39:0] _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1_string;
  reg [39:0] _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2_string;
  reg [31:0] _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_string;
  reg [31:0] _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_1_string;
  reg [31:0] _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_2_string;
  reg [79:0] _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1_string;
  reg [79:0] _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_string;
  reg [79:0] _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_3_string;
  reg [79:0] LsuPlugin_logic_flusher_stateReg_string;
  reg [79:0] LsuPlugin_logic_flusher_stateNext_string;
  reg [87:0] TrapPlugin_logic_harts_0_trap_fsm_stateReg_string;
  reg [87:0] TrapPlugin_logic_harts_0_trap_fsm_stateNext_string;
  reg [47:0] MmuPlugin_logic_refill_stateReg_string;
  reg [47:0] MmuPlugin_logic_refill_stateNext_string;
  reg [71:0] PerformanceCounterPlugin_logic_fsm_stateReg_string;
  reg [71:0] PerformanceCounterPlugin_logic_fsm_stateNext_string;
  reg [79:0] CsrAccessPlugin_logic_fsm_stateReg_string;
  reg [79:0] CsrAccessPlugin_logic_fsm_stateNext_string;
  `endif

  (* ram_style = "distributed" *) reg [37:0] BtbPlugin_logic_ras_mem_stack [0:3];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol0 [0:511];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol1 [0:511];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol2 [0:511];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol3 [0:511];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol4 [0:511];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol5 [0:511];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol6 [0:511];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol7 [0:511];
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_1;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_2;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_3;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_4;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_5;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_6;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_7;
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol0 [0:511];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol1 [0:511];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol2 [0:511];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol3 [0:511];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol4 [0:511];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol5 [0:511];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol6 [0:511];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol7 [0:511];
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_1;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_2;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_3;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_4;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_5;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_6;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_7;
  reg [21:0] LsuL1Plugin_logic_ways_0_mem [0:63];
  reg [21:0] LsuL1Plugin_logic_ways_1_mem [0:63];
  reg [2:0] LsuL1Plugin_logic_shared_mem [0:63];
  reg [63:0] LsuL1Plugin_logic_writeback_victimBuffer [0:7];
  reg [63:0] FetchL1Plugin_logic_banks_0_mem [0:511];
  reg [63:0] FetchL1Plugin_logic_banks_1_mem [0:511];
  reg [21:0] FetchL1Plugin_logic_ways_0_mem [0:63];
  reg [21:0] FetchL1Plugin_logic_ways_1_mem [0:63];
  reg [0:0] FetchL1Plugin_logic_plru_mem [0:63];
  reg [3:0] GSharePlugin_logic_mem_banks_0 [0:8191];
  (* ram_style = "block" *) reg [57:0] BtbPlugin_logic_mem [0:511];
  (* ram_style = "distributed" *) reg [46:0] FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_0 [0:31];
  (* ram_style = "distributed" *) reg [46:0] FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_1 [0:31];
  (* ram_style = "distributed" *) reg [28:0] FetchL1Plugin_logic_translationStorage_logic_sl_1_ways_0 [0:31];
  (* ram_style = "distributed" *) reg [46:0] LsuPlugin_logic_translationStorage_logic_sl_0_ways_0 [0:31];
  (* ram_style = "distributed" *) reg [46:0] LsuPlugin_logic_translationStorage_logic_sl_0_ways_1 [0:31];
  (* ram_style = "distributed" *) reg [46:0] LsuPlugin_logic_translationStorage_logic_sl_0_ways_2 [0:31];
  (* ram_style = "distributed" *) reg [28:0] LsuPlugin_logic_translationStorage_logic_sl_1_ways_0 [0:31];
  reg [63:0] CsrRamPlugin_logic_mem [0:15];
  function [2:0] zz_FetchL1Plugin_logic_trapPort_payload_arg(input dummy);
    begin
      zz_FetchL1Plugin_logic_trapPort_payload_arg = 3'b000;
      zz_FetchL1Plugin_logic_trapPort_payload_arg[1 : 0] = 2'b10;
      zz_FetchL1Plugin_logic_trapPort_payload_arg[2 : 2] = 1'b0;
    end
  endfunction
  wire [2:0] _zz_60;

  assign _zz_when_1 = (! FetchL1Plugin_logic_refill_slots_0_valid);
  assign _zz_PmpPlugin_logic_entries_0_napot_24 = ({1'd0,_zz_PmpPlugin_logic_entries_0_napot_16} <<< 1'd1);
  assign _zz_PmpPlugin_logic_entries_1_napot_24 = ({1'd0,_zz_PmpPlugin_logic_entries_1_napot_16} <<< 1'd1);
  assign _zz_PmpPlugin_logic_entries_2_napot_24 = ({1'd0,_zz_PmpPlugin_logic_entries_2_napot_16} <<< 1'd1);
  assign _zz_PmpPlugin_logic_entries_3_napot_24 = ({1'd0,_zz_PmpPlugin_logic_entries_3_napot_16} <<< 1'd1);
  assign _zz_early0_IntAluPlugin_logic_alu_result = (early0_IntAluPlugin_logic_alu_bitwise | _zz_early0_IntAluPlugin_logic_alu_result_1);
  assign _zz_early0_IntAluPlugin_logic_alu_result_1 = (execute_ctrl2_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0 ? execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0 : 64'h0);
  assign _zz_early0_IntAluPlugin_logic_alu_result_2 = (execute_ctrl2_down_early0_IntAluPlugin_ALU_SLTX_lane0 ? _zz_early0_IntAluPlugin_logic_alu_result_3 : 64'h0);
  assign _zz_early0_IntAluPlugin_logic_alu_result_3 = _zz_early0_IntAluPlugin_logic_alu_result_4;
  assign _zz_early0_IntAluPlugin_logic_alu_result_5 = execute_ctrl2_down_early0_SrcPlugin_LESS_lane0;
  assign _zz_early0_IntAluPlugin_logic_alu_result_4 = {63'd0, _zz_early0_IntAluPlugin_logic_alu_result_5};
  assign _zz_early0_BarrelShifterPlugin_logic_shift_amplitude = execute_ctrl2_down_early0_SrcPlugin_SRC2_lane0[5 : 0];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_reversed = {execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[0],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[1],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[2],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[3],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[4],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[5],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[6],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[7],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[8],{_zz_early0_BarrelShifterPlugin_logic_shift_reversed_1,{_zz_early0_BarrelShifterPlugin_logic_shift_reversed_2,_zz_early0_BarrelShifterPlugin_logic_shift_reversed_3}}}}}}}}}}};
  assign _zz_early0_BarrelShifterPlugin_logic_shift_shifted = ($signed(_zz_early0_BarrelShifterPlugin_logic_shift_shifted_1) >>> early0_BarrelShifterPlugin_logic_shift_amplitude);
  assign _zz_early0_BarrelShifterPlugin_logic_shift_shifted_1 = {(execute_ctrl2_down_BarrelShifterPlugin_SIGNED_lane0 && execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[63]),early0_BarrelShifterPlugin_logic_shift_reversed};
  assign _zz_early0_BarrelShifterPlugin_logic_shift_patched = {early0_BarrelShifterPlugin_logic_shift_shifted[0],{early0_BarrelShifterPlugin_logic_shift_shifted[1],{early0_BarrelShifterPlugin_logic_shift_shifted[2],{early0_BarrelShifterPlugin_logic_shift_shifted[3],{early0_BarrelShifterPlugin_logic_shift_shifted[4],{early0_BarrelShifterPlugin_logic_shift_shifted[5],{early0_BarrelShifterPlugin_logic_shift_shifted[6],{early0_BarrelShifterPlugin_logic_shift_shifted[7],{early0_BarrelShifterPlugin_logic_shift_shifted[8],{_zz_early0_BarrelShifterPlugin_logic_shift_patched_1,{_zz_early0_BarrelShifterPlugin_logic_shift_patched_2,_zz_early0_BarrelShifterPlugin_logic_shift_patched_3}}}}}}}}}}};
  assign _zz_LsuL1Plugin_logic_shared_lsuRead_rsp_plru_0_1 = _zz_LsuL1Plugin_logic_shared_lsuRead_rsp_plru_0[0 : 0];
  assign _zz_LsuL1Plugin_logic_writeback_read_wordIndex_1 = LsuL1Plugin_logic_writeback_read_slotRead_valid;
  assign _zz_LsuL1Plugin_logic_writeback_read_wordIndex = {2'd0, _zz_LsuL1Plugin_logic_writeback_read_wordIndex_1};
  assign _zz_LsuL1Plugin_logic_writeback_write_wordIndex_1 = (LsuL1Plugin_logic_writeback_write_bufferRead_fire && 1'b1);
  assign _zz_LsuL1Plugin_logic_writeback_write_wordIndex = {2'd0, _zz_LsuL1Plugin_logic_writeback_write_wordIndex_1};
  assign _zz_LsuL1Plugin_logic_lsu_ctrl_refillWayNeedWriteback = ({execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_loaded,execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_loaded} & execute_ctrl4_down_LsuL1Plugin_logic_SHARED_lane0_dirty);
  assign _zz_LsuL1Plugin_logic_lsu_ctrl_doWrite = ((_zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0 ? (1'b1 && (! execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault)) : 1'b0) | (_zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0_1 ? (1'b1 && (! execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault)) : 1'b0));
  assign _zz_LsuL1Plugin_logic_shared_write_payload_data_dirty = (2'b01 <<< LsuL1Plugin_logic_lsu_ctrl_refillWayWithoutUpdate);
  assign _zz_when = 1'b1;
  assign _zz_LsuL1Plugin_logic_waysWrite_tag_fault = ((_zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0 ? execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault : 1'b0) | (_zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0_1 ? execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault : 1'b0));
  assign _zz_LsuL1Plugin_logic_shared_write_payload_data_plru_0_1 = _zz_LsuL1Plugin_logic_shared_write_payload_data_plru_0[0 : 0];
  assign _zz_execute_ctrl2_down_MUL_SRC1_lane0 = {(execute_ctrl2_down_RsUnsignedPlugin_RS1_SIGNED_lane0 && execute_ctrl2_up_integer_RS1_lane0[63]),execute_ctrl2_up_integer_RS1_lane0};
  assign _zz_execute_ctrl2_down_MUL_SRC2_lane0 = {(execute_ctrl2_down_RsUnsignedPlugin_RS2_SIGNED_lane0 && execute_ctrl2_up_integer_RS2_lane0[63]),execute_ctrl2_up_integer_RS2_lane0};
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_6_lane0_1 = ($signed(_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_6_lane0_2) * $signed(_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_6_lane0_3));
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_6_lane0 = {{45{_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_6_lane0_1[31]}}, _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_6_lane0_1};
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_6_lane0_2 = {1'b0,execute_ctrl2_down_MUL_SRC1_lane0[16 : 0]};
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_6_lane0_3 = execute_ctrl2_down_MUL_SRC2_lane0[64 : 51];
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_7_lane0_1 = ($signed(_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_7_lane0_2) * $signed(_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_7_lane0_3));
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_7_lane0 = {{45{_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_7_lane0_1[31]}}, _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_7_lane0_1};
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_7_lane0_2 = execute_ctrl2_down_MUL_SRC1_lane0[64 : 51];
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_7_lane0_3 = {1'b0,execute_ctrl2_down_MUL_SRC2_lane0[16 : 0]};
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_10_lane0_1 = ($signed(_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_10_lane0_2) * $signed(_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_10_lane0_3));
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_10_lane0 = {{28{_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_10_lane0_1[31]}}, _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_10_lane0_1};
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_10_lane0_2 = {1'b0,execute_ctrl2_down_MUL_SRC1_lane0[33 : 17]};
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_10_lane0_3 = execute_ctrl2_down_MUL_SRC2_lane0[64 : 51];
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_11_lane0_1 = ($signed(_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_11_lane0_2) * $signed(_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_11_lane0_3));
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_11_lane0 = {{28{_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_11_lane0_1[31]}}, _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_11_lane0_1};
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_11_lane0_2 = execute_ctrl2_down_MUL_SRC1_lane0[64 : 51];
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_11_lane0_3 = {1'b0,execute_ctrl2_down_MUL_SRC2_lane0[33 : 17]};
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_13_lane0_1 = ($signed(_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_13_lane0_2) * $signed(_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_13_lane0_3));
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_13_lane0 = {{11{_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_13_lane0_1[31]}}, _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_13_lane0_1};
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_13_lane0_2 = {1'b0,execute_ctrl2_down_MUL_SRC1_lane0[50 : 34]};
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_13_lane0_3 = execute_ctrl2_down_MUL_SRC2_lane0[64 : 51];
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_14_lane0_1 = ($signed(_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_14_lane0_2) * $signed(_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_14_lane0_3));
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_14_lane0 = {{11{_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_14_lane0_1[31]}}, _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_14_lane0_1};
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_14_lane0_2 = execute_ctrl2_down_MUL_SRC1_lane0[64 : 51];
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_14_lane0_3 = {1'b0,execute_ctrl2_down_MUL_SRC2_lane0[50 : 34]};
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_15_lane0_1 = ($signed(_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_15_lane0_2) * $signed(_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_15_lane0_3));
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_15_lane0 = _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_15_lane0_1[25:0];
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_15_lane0_2 = execute_ctrl2_down_MUL_SRC1_lane0[64 : 51];
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_15_lane0_3 = execute_ctrl2_down_MUL_SRC2_lane0[64 : 51];
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_7 = (_zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_8 + _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_11);
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_8 = (_zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_9 + _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_10);
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_9 = {3'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_10 = {3'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_1};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_11 = (_zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_12 + _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_13);
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_12 = {3'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_2};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_13 = {3'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_3};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_14 = (_zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_15 + _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_18);
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_15 = (_zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_16 + _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_17);
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_16 = {3'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_4};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_17 = {3'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_5};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_18 = {3'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_6};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_7 = (_zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_8 + _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_11);
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_8 = (_zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_9 + _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_10);
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_9 = {3'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_10 = {3'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_1};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_11 = (_zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_12 + _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_13);
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_12 = {3'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_2};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_13 = {3'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_3};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_14 = (_zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_15 + _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_18);
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_15 = (_zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_16 + _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_17);
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_16 = {3'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_4};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_17 = {3'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_5};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_18 = {3'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_6};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_7 = (_zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_8 + _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_11);
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_8 = (_zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_9 + _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_10);
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_9 = {3'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_10 = {3'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_1};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_11 = (_zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_12 + _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_13);
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_12 = {3'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_2};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_13 = {3'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_3};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_14 = (_zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_15 + _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_18);
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_15 = (_zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_16 + _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_17);
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_16 = {3'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_4};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_17 = {3'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_5};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_18 = {3'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_6};
  assign _zz_execute_ctrl2_down_RsUnsignedPlugin_RS1_UNSIGNED_lane0_1 = execute_ctrl2_down_RsUnsignedPlugin_RS1_REVERT_lane0;
  assign _zz_execute_ctrl2_down_RsUnsignedPlugin_RS1_UNSIGNED_lane0 = {63'd0, _zz_execute_ctrl2_down_RsUnsignedPlugin_RS1_UNSIGNED_lane0_1};
  assign _zz_execute_ctrl2_down_RsUnsignedPlugin_RS2_UNSIGNED_lane0_1 = execute_ctrl2_down_RsUnsignedPlugin_RS2_REVERT_lane0;
  assign _zz_execute_ctrl2_down_RsUnsignedPlugin_RS2_UNSIGNED_lane0 = {63'd0, _zz_execute_ctrl2_down_RsUnsignedPlugin_RS2_UNSIGNED_lane0_1};
  assign _zz_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0_1 = ((early0_DivPlugin_logic_processing_divRevertResult ? (~ _zz_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0) : _zz_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0) + _zz_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0_2);
  assign _zz_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0_3 = early0_DivPlugin_logic_processing_divRevertResult;
  assign _zz_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0_2 = {63'd0, _zz_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0_3};
  assign _zz_FetchL1Plugin_logic_hits_w_0_indirect_bypassHits = {7'd0, fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_address};
  assign _zz_FetchL1Plugin_logic_hits_w_0_indirect_bypassHits_1 = (fetch_logic_ctrls_1_down_Fetch_WORD_PC >>> 4'd12);
  assign _zz_FetchL1Plugin_logic_hits_w_1_indirect_bypassHits = {7'd0, fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_address};
  assign _zz_FetchL1Plugin_logic_hits_w_1_indirect_bypassHits_1 = (fetch_logic_ctrls_1_down_Fetch_WORD_PC >>> 4'd12);
  assign _zz_FetchL1Plugin_logic_ctrl_dataAccessFault = ((fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_0 ? fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_0_error : 1'b0) | (fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_1 ? fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_1_error : 1'b0));
  assign _zz_FetchL1Plugin_logic_plru_write_payload_data_0 = 1'b0;
  assign _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_5 = fetch_logic_ctrls_0_down_Prediction_BRANCH_HISTORY;
  assign _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_4 = {1'd0, _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_5};
  assign _zz_BtbPlugin_logic_ras_ptr_push = (BtbPlugin_logic_ras_ptr_push + _zz_BtbPlugin_logic_ras_ptr_push_1);
  assign _zz_BtbPlugin_logic_ras_ptr_push_2 = BtbPlugin_logic_ras_ptr_pushIt;
  assign _zz_BtbPlugin_logic_ras_ptr_push_1 = {1'd0, _zz_BtbPlugin_logic_ras_ptr_push_2};
  assign _zz_BtbPlugin_logic_ras_ptr_push_4 = BtbPlugin_logic_ras_ptr_popIt;
  assign _zz_BtbPlugin_logic_ras_ptr_push_3 = {1'd0, _zz_BtbPlugin_logic_ras_ptr_push_4};
  assign _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue = (BtbPlugin_logic_ras_ptr_pop + _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_1);
  assign _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_2 = BtbPlugin_logic_ras_ptr_pushIt;
  assign _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_1 = {1'd0, _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_2};
  assign _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_4 = BtbPlugin_logic_ras_ptr_popIt;
  assign _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_3 = {1'd0, _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_4};
  assign _zz_WhiteboxerPlugin_logic_decodes_0_pc_1 = decode_ctrls_0_down_PC_0;
  assign _zz_WhiteboxerPlugin_logic_decodes_0_pc = {{25{_zz_WhiteboxerPlugin_logic_decodes_0_pc_1[38]}}, _zz_WhiteboxerPlugin_logic_decodes_0_pc_1};
  assign _zz_FetchL1Plugin_pmaBuilder_onTransfers_0_addressHit = (|_zz_FetchL1Plugin_logic_ctrl_pmaPort_rsp_io);
  assign _zz_FetchL1Plugin_logic_ctrl_pmaPort_rsp_io_1 = (|_zz_FetchL1Plugin_logic_ctrl_pmaPort_rsp_io);
  assign _zz_PerformanceCounterPlugin_logic_eventInstructions_0 = ((! PerformanceCounterPlugin_logic_ignoreNextCommit) ? PerformanceCounterPlugin_logic_commitMask : 1'b0);
  assign _zz_PerformanceCounterPlugin_logic_counters_cycle_value_1 = (! PerformanceCounterPlugin_logic_counters_cycle_mcountinhibit);
  assign _zz_PerformanceCounterPlugin_logic_counters_cycle_value = {7'd0, _zz_PerformanceCounterPlugin_logic_counters_cycle_value_1};
  assign _zz_PerformanceCounterPlugin_logic_counters_instret_value_1 = {7'd0, _zz_PerformanceCounterPlugin_logic_counters_instret_value};
  assign _zz_LsuPlugin_logic_onAddress0_ls_port_payload_address = execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0;
  assign _zz_LsuPlugin_logic_onAddress0_ls_storeId_1 = LsuPlugin_logic_onAddress0_ls_port_fire;
  assign _zz_LsuPlugin_logic_onAddress0_ls_storeId = {11'd0, _zz_LsuPlugin_logic_onAddress0_ls_storeId_1};
  assign _zz_LsuPlugin_logic_onAddress0_flush_port_payload_address = ({6'd0,LsuPlugin_logic_flusher_cmdCounter} <<< 3'd6);
  assign _zz_LsuPlugin_logic_onPma_addressExtension = execute_ctrl3_down_early0_SrcPlugin_ADD_SUB_lane0;
  assign _zz__zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0 = execute_ctrl3_down_early0_SrcPlugin_ADD_SUB_lane0[63 : 39];
  assign _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub = ($signed(_zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_1) + $signed(_zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_4));
  assign _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_1 = ($signed(_zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_2) + $signed(_zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_3));
  assign _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_2 = execute_ctrl4_up_integer_RS2_lane0;
  assign _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_3 = (LsuPlugin_logic_onCtrl_rva_alu_compare ? (~ LsuPlugin_logic_onCtrl_rva_srcBuffer) : LsuPlugin_logic_onCtrl_rva_srcBuffer);
  assign _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_5 = (LsuPlugin_logic_onCtrl_rva_alu_compare ? 2'b01 : 2'b00);
  assign _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_4 = {{62{_zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_5[1]}}, _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_5};
  assign _zz_LsuPlugin_logic_trapPort_payload_code = (execute_ctrl4_down_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0 ? (execute_ctrl4_down_LsuL1_STORE_lane0 ? 3'b110 : 3'b100) : 3'b000);
  assign _zz_LsuPlugin_logic_flusher_cmdCounter = execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0[11 : 6];
  assign _zz__zz_execute_ctrl1_down_early0_SrcPlugin_SRC1_lane0 = {execute_ctrl1_down_Decode_UOP_lane0[31 : 12],12'h0};
  assign _zz__zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0 = execute_ctrl1_down_Decode_UOP_lane0[31 : 20];
  assign _zz__zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0_1 = execute_ctrl1_down_PC_lane0;
  assign _zz__zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0_2 = {execute_ctrl1_down_Decode_UOP_lane0[31 : 25],execute_ctrl1_down_Decode_UOP_lane0[11 : 7]};
  assign _zz_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0 = ($signed(execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0) + $signed(early0_SrcPlugin_logic_addsub_combined_rs2Patched));
  assign _zz_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0_1 = _zz_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0_2;
  assign _zz_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0_3 = execute_ctrl2_down_SrcStageables_REVERT_lane0;
  assign _zz_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0_2 = {63'd0, _zz_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0_3};
  assign _zz_early0_BranchPlugin_pcCalc_target_b = {{{{execute_ctrl2_down_Decode_UOP_lane0[31],execute_ctrl2_down_Decode_UOP_lane0[19 : 12]},execute_ctrl2_down_Decode_UOP_lane0[20]},execute_ctrl2_down_Decode_UOP_lane0[30 : 21]},1'b0};
  assign _zz_early0_BranchPlugin_pcCalc_target_b_1 = execute_ctrl2_down_Decode_UOP_lane0[31 : 20];
  assign _zz_early0_BranchPlugin_pcCalc_target_b_2 = {{{{execute_ctrl2_down_Decode_UOP_lane0[31],execute_ctrl2_down_Decode_UOP_lane0[7]},execute_ctrl2_down_Decode_UOP_lane0[30 : 25]},execute_ctrl2_down_Decode_UOP_lane0[11 : 8]},1'b0};
  assign _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0 = _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0_1;
  assign _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0_1 = ($signed(_zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0_2) + $signed(early0_BranchPlugin_pcCalc_target_b));
  assign _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0_2 = {{25{early0_BranchPlugin_pcCalc_target_a[38]}}, early0_BranchPlugin_pcCalc_target_a};
  assign _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0_1 = ({1'd0,early0_BranchPlugin_pcCalc_slices} <<< 1'd1);
  assign _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0 = {36'd0, _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0_1};
  assign _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0_1 = ({1'd0,execute_ctrl2_down_Decode_INSTRUCTION_SLICE_COUNT_lane0} <<< 1'd1);
  assign _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0 = {37'd0, _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0_1};
  assign _zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_LAST = (2'b01 <<< fetch_logic_ctrls_2_down_Prediction_WORD_JUMP_SLICE);
  assign _zz_AlignerPlugin_logic_extractors_0_redo_4 = (((_zz_AlignerPlugin_logic_extractors_0_redo ? AlignerPlugin_logic_scanners_0_redo : 1'b0) | (_zz_AlignerPlugin_logic_extractors_0_redo_1 ? AlignerPlugin_logic_scanners_1_redo : 1'b0)) | ((_zz_AlignerPlugin_logic_extractors_0_redo_2 ? AlignerPlugin_logic_scanners_2_redo : 1'b0) | (_zz_AlignerPlugin_logic_extractors_0_redo_3 ? AlignerPlugin_logic_scanners_3_redo : 1'b0)));
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_22 = {{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_7,AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 2]},12'h0};
  assign _zz__zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_18_1 = {AlignerPlugin_logic_extractors_0_ctx_instruction[12],AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 2]};
  assign _zz__zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_18 = {6'd0, _zz__zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_18_1};
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_31 = {{{4'b0000,AlignerPlugin_logic_extractors_0_ctx_instruction[8 : 7]},AlignerPlugin_logic_extractors_0_ctx_instruction[12 : 9]},2'b00};
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_32 = {{{4'b0000,AlignerPlugin_logic_extractors_0_ctx_instruction[8 : 7]},AlignerPlugin_logic_extractors_0_ctx_instruction[12 : 9]},2'b00};
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_33 = {{{3'b000,AlignerPlugin_logic_extractors_0_ctx_instruction[9 : 7]},AlignerPlugin_logic_extractors_0_ctx_instruction[12 : 10]},3'b000};
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_34 = {{{3'b000,AlignerPlugin_logic_extractors_0_ctx_instruction[9 : 7]},AlignerPlugin_logic_extractors_0_ctx_instruction[12 : 10]},3'b000};
  assign _zz__zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_5 = {_zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_4[0],_zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_4[1]};
  assign _zz_early0_EnvPlugin_logic_trapPort_payload_tval_1 = ((|{(execute_ctrl2_down_early0_EnvPlugin_OP_lane0 == EnvPluginOp_SFENCE_VMA),{(execute_ctrl2_down_early0_EnvPlugin_OP_lane0 == EnvPluginOp_WFI),(execute_ctrl2_down_early0_EnvPlugin_OP_lane0 == EnvPluginOp_PRIV_RET)}}) ? execute_ctrl2_down_Decode_UOP_lane0 : 32'h0);
  assign _zz_early0_EnvPlugin_logic_trapPort_payload_tval = {7'd0, _zz_early0_EnvPlugin_logic_trapPort_payload_tval_1};
  assign _zz_early0_EnvPlugin_logic_trapPort_payload_code = {2'd0, early0_EnvPlugin_logic_exe_privilege};
  assign _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_napot_MATCH = ({12'd0,PmpPlugin_logic_entries_0_address[20 : 1]} <<< 4'd12);
  assign _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_tor_BIGGER = (PmpPlugin_logic_entries_0_address >>> 1'd1);
  assign _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_napot_MATCH = ({12'd0,PmpPlugin_logic_entries_1_address[20 : 1]} <<< 4'd12);
  assign _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_tor_BIGGER = (PmpPlugin_logic_entries_1_address >>> 1'd1);
  assign _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_napot_MATCH = ({12'd0,PmpPlugin_logic_entries_2_address[20 : 1]} <<< 4'd12);
  assign _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_tor_BIGGER = (PmpPlugin_logic_entries_2_address >>> 1'd1);
  assign _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_napot_MATCH = ({12'd0,PmpPlugin_logic_entries_3_address[20 : 1]} <<< 4'd12);
  assign _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_tor_BIGGER = (PmpPlugin_logic_entries_3_address >>> 1'd1);
  assign _zz_fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_ACCESS_FAULT_4 = (((_zz_fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_ACCESS_FAULT ? PmpPlugin_logic_entries_0_isLocked : 1'b0) | (_zz_fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_ACCESS_FAULT_1 ? PmpPlugin_logic_entries_1_isLocked : 1'b0)) | ((_zz_fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_ACCESS_FAULT_2 ? PmpPlugin_logic_entries_2_isLocked : 1'b0) | (_zz_fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_ACCESS_FAULT_3 ? PmpPlugin_logic_entries_3_isLocked : 1'b0)));
  assign _zz_fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_ACCESS_FAULT_5 = (((_zz_fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_ACCESS_FAULT ? fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_PERM_OK : 1'b0) | (_zz_fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_ACCESS_FAULT_1 ? fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_PERM_OK : 1'b0)) | ((_zz_fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_ACCESS_FAULT_2 ? fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_PERM_OK : 1'b0) | (_zz_fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_ACCESS_FAULT_3 ? fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_PERM_OK : 1'b0)));
  assign _zz_execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_0_napot_MATCH_lane0 = ({12'd0,PmpPlugin_logic_entries_0_address[20 : 1]} <<< 4'd12);
  assign _zz_execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_0_tor_BIGGER_lane0 = (PmpPlugin_logic_entries_0_address >>> 1'd1);
  assign _zz_execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_1_napot_MATCH_lane0 = ({12'd0,PmpPlugin_logic_entries_1_address[20 : 1]} <<< 4'd12);
  assign _zz_execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_1_tor_BIGGER_lane0 = (PmpPlugin_logic_entries_1_address >>> 1'd1);
  assign _zz_execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_2_napot_MATCH_lane0 = ({12'd0,PmpPlugin_logic_entries_2_address[20 : 1]} <<< 4'd12);
  assign _zz_execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_2_tor_BIGGER_lane0 = (PmpPlugin_logic_entries_2_address >>> 1'd1);
  assign _zz_execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_3_napot_MATCH_lane0 = ({12'd0,PmpPlugin_logic_entries_3_address[20 : 1]} <<< 4'd12);
  assign _zz_execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_3_tor_BIGGER_lane0 = (PmpPlugin_logic_entries_3_address >>> 1'd1);
  assign _zz_execute_ctrl4_down_LsuPlugin_logic_pmpPort_ACCESS_FAULT_lane0_4 = (((_zz_execute_ctrl4_down_LsuPlugin_logic_pmpPort_ACCESS_FAULT_lane0 ? PmpPlugin_logic_entries_0_isLocked : 1'b0) | (_zz_execute_ctrl4_down_LsuPlugin_logic_pmpPort_ACCESS_FAULT_lane0_1 ? PmpPlugin_logic_entries_1_isLocked : 1'b0)) | ((_zz_execute_ctrl4_down_LsuPlugin_logic_pmpPort_ACCESS_FAULT_lane0_2 ? PmpPlugin_logic_entries_2_isLocked : 1'b0) | (_zz_execute_ctrl4_down_LsuPlugin_logic_pmpPort_ACCESS_FAULT_lane0_3 ? PmpPlugin_logic_entries_3_isLocked : 1'b0)));
  assign _zz_execute_ctrl4_down_LsuPlugin_logic_pmpPort_ACCESS_FAULT_lane0_5 = (((_zz_execute_ctrl4_down_LsuPlugin_logic_pmpPort_ACCESS_FAULT_lane0 ? execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_0_PERM_OK_lane0 : 1'b0) | (_zz_execute_ctrl4_down_LsuPlugin_logic_pmpPort_ACCESS_FAULT_lane0_1 ? execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_1_PERM_OK_lane0 : 1'b0)) | ((_zz_execute_ctrl4_down_LsuPlugin_logic_pmpPort_ACCESS_FAULT_lane0_2 ? execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_2_PERM_OK_lane0 : 1'b0) | (_zz_execute_ctrl4_down_LsuPlugin_logic_pmpPort_ACCESS_FAULT_lane0_3 ? execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_3_PERM_OK_lane0 : 1'b0)));
  assign _zz_LsuPlugin_pmaBuilder_l1_onTransfers_0_addressHit = (|_zz_LsuPlugin_logic_onPma_cached_rsp_io);
  assign _zz_LsuPlugin_logic_onPma_cached_rsp_io_1 = (|_zz_LsuPlugin_logic_onPma_cached_rsp_io);
  assign _zz_LsuPlugin_pmaBuilder_io_onTransfers_0_addressHit = (|((LsuPlugin_pmaBuilder_io_addressBits & 32'h0) == 32'h0));
  assign _zz_LsuPlugin_logic_onPma_io_rsp_io = (|((LsuPlugin_pmaBuilder_io_addressBits & 32'h70000000) == 32'h0));
  assign _zz_early0_BranchPlugin_logic_alu_expectedMsb = execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0;
  assign _zz__zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0 = execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[63 : 39];
  assign _zz_early0_BranchPlugin_logic_jumpLogic_history_shifter_1 = {early0_BranchPlugin_logic_jumpLogic_history_shifter,execute_ctrl2_down_Prediction_ALIGNED_SLICES_TAKEN_lane0[0]};
  assign _zz_early0_BranchPlugin_logic_jumpLogic_history_shifter_2 = {early0_BranchPlugin_logic_jumpLogic_history_shifter_1,execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0};
  assign _zz_early0_BranchPlugin_logic_wb_payload_1 = execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0;
  assign _zz_early0_BranchPlugin_logic_wb_payload = {{25{_zz_early0_BranchPlugin_logic_wb_payload_1[38]}}, _zz_early0_BranchPlugin_logic_wb_payload_1};
  assign _zz_decode_ctrls_1_down_RS1_ENABLE_0 = (|{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000044) == 32'h0),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000018) == 32'h0),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00006004) == 32'h00002000),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & _zz_decode_ctrls_1_down_RS1_ENABLE_0_1) == 32'h00001000),((decode_ctrls_1_down_Decode_INSTRUCTION_0 & _zz_decode_ctrls_1_down_RS1_ENABLE_0_2) == 32'h00002000)}}}});
  assign _zz_decode_ctrls_1_down_RS1_PHYS_0 = decode_ctrls_1_down_Decode_INSTRUCTION_0[19 : 15];
  assign _zz_decode_ctrls_1_down_RS2_ENABLE_0 = (|{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000034) == 32'h00000020),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000064) == 32'h00000020),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h08000070) == 32'h08000020),((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h10000070) == 32'h00000020)}}});
  assign _zz_decode_ctrls_1_down_RS2_PHYS_0 = decode_ctrls_1_down_Decode_INSTRUCTION_0[24 : 20];
  assign _zz_decode_ctrls_1_down_RD_ENABLE_0 = (|{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000028) == 32'h00000028),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00001010) == 32'h00001010),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00002010) == 32'h00002010),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & _zz_decode_ctrls_1_down_RD_ENABLE_0_1) == 32'h00000010),{(_zz_decode_ctrls_1_down_RD_ENABLE_0_2 == _zz_decode_ctrls_1_down_RD_ENABLE_0_3),(_zz_decode_ctrls_1_down_RD_ENABLE_0_4 == _zz_decode_ctrls_1_down_RD_ENABLE_0_5)}}}}});
  assign _zz_decode_ctrls_1_down_RD_PHYS_0 = decode_ctrls_1_down_Decode_INSTRUCTION_0[11 : 7];
  assign _zz_DecoderPlugin_logic_laneLogic_0_fixer_isJb = (|((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000050) == 32'h00000040));
  assign _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice_1 = ((! decode_ctrls_1_down_Prediction_ALIGN_REDO_0) ? _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice_2 : 2'b00);
  assign _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice = {37'd0, _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice_1};
  assign _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice_2 = ({1'd0,decode_ctrls_1_down_Decode_INSTRUCTION_SLICE_COUNT_0} <<< 1'd1);
  assign _zz_GSharePlugin_logic_onLearn_hash_5 = LearnPlugin_logic_learn_payload_history;
  assign _zz_GSharePlugin_logic_onLearn_hash_4 = {1'd0, _zz_GSharePlugin_logic_onLearn_hash_5};
  assign _zz_BtbPlugin_logic_memWrite_payload_address = (LearnPlugin_logic_learn_payload_pcOnLastSlice >>> 2'd2);
  assign _zz_decode_ctrls_1_down_AguPlugin_CLEAN_0 = _zz_decode_ctrls_1_down_AguPlugin_CLEAN_0_1[0];
  assign _zz_decode_ctrls_1_down_AguPlugin_CLEAN_0_1 = (|{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00102028) == 32'h00102008),((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00202028) == 32'h00202008)});
  assign _zz_decode_ctrls_1_down_AguPlugin_INVALIDATE_0 = _zz_decode_ctrls_1_down_AguPlugin_INVALIDATE_0_1[0];
  assign _zz_decode_ctrls_1_down_AguPlugin_INVALIDATE_0_1 = (|((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00302028) == 32'h00002008));
  assign _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_0 = _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_0_1[0];
  assign _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_0_1 = 1'b0;
  assign _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_0 = _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_0_1[0];
  assign _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_0_1 = 1'b0;
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0_1[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0_1 = (|_zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_0 = _zz_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_0_1[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_0_1 = (|{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000040) == 32'h00000040),((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000010) == 32'h0)});
  assign _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_0 = _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_0_1[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_0_1 = (|{_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_1,_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0});
  assign _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_0 = _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_0_1[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_0_1 = (|{_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_1,_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0});
  assign _zz_decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_0 = _zz_decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_0_1[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_0_1 = (|{_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_1,_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0});
  assign _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_0 = _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_0_1[0];
  assign _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_0_1 = (|{_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_1,_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0});
  assign _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_2 = _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_3[0];
  assign _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_3 = (|{_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_1,_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0});
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_0 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_0_1[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_0_1 = (|_zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0_1 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0_2[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0_2 = (|_zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0);
  assign _zz_BtbPlugin_logic_memWrite_payload_address_1 = (DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice >>> 2'd2);
  assign _zz_BtbPlugin_logic_memRead_cmd_payload = (fetch_logic_ctrls_0_down_Fetch_WORD_PC >>> 2'd2);
  assign _zz_BtbPlugin_logic_ras_write_payload_data = (BtbPlugin_logic_applyIt_rasLogic_pushPc + 39'h0000000002);
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_slices = {1'd0, execute_ctrl4_down_Decode_INSTRUCTION_SLICE_COUNT_lane0};
  assign _zz_TrapPlugin_logic_harts_0_trap_fsm_jumpTarget_1 = ({1'd0,TrapPlugin_logic_harts_0_trap_fsm_jumpOffset} <<< 1'd1);
  assign _zz_TrapPlugin_logic_harts_0_trap_fsm_jumpTarget = {36'd0, _zz_TrapPlugin_logic_harts_0_trap_fsm_jumpTarget_1};
  assign _zz_PcPlugin_logic_harts_0_self_pc_1 = (PcPlugin_logic_harts_0_self_increment ? 3'b100 : 3'b000);
  assign _zz_PcPlugin_logic_harts_0_self_pc = {36'd0, _zz_PcPlugin_logic_harts_0_self_pc_1};
  assign _zz_PcPlugin_logic_harts_0_aggregator_fault = (((_zz_PcPlugin_logic_harts_0_aggregator_target ? TrapPlugin_logic_harts_0_trap_pcPort_payload_fault : 1'b0) | (_zz_PcPlugin_logic_harts_0_aggregator_target_1 ? early0_BranchPlugin_logic_pcPort_payload_fault : 1'b0)) | (_zz_PcPlugin_logic_harts_0_aggregator_target_2 ? PcPlugin_logic_harts_0_self_flow_payload_fault : 1'b0));
  assign _zz_PcPlugin_logic_harts_0_aggregator_fault_1_1 = (_zz_PcPlugin_logic_harts_0_aggregator_fault_1 ? BtbPlugin_logic_pcPort_payload_fault : 1'b0);
  assign _zz_LsuPlugin_logic_translationStorage_logic_sl_0_allocId_valueNext_1 = LsuPlugin_logic_translationStorage_logic_sl_0_allocId_willIncrement;
  assign _zz_LsuPlugin_logic_translationStorage_logic_sl_0_allocId_valueNext = {1'd0, _zz_LsuPlugin_logic_translationStorage_logic_sl_0_allocId_valueNext_1};
  assign _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_4 = (((_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute ? execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_allowExecute : 1'b0) | (_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_1 ? execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_allowExecute : 1'b0)) | ((_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_2 ? execute_ctrl3_down_MMU_L0_ENTRIES_lane0_2_allowExecute : 1'b0) | (_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_3 ? execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_allowExecute : 1'b0)));
  assign _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowRead = (((_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute ? execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_allowRead : 1'b0) | (_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_1 ? execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_allowRead : 1'b0)) | ((_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_2 ? execute_ctrl3_down_MMU_L0_ENTRIES_lane0_2_allowRead : 1'b0) | (_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_3 ? execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_allowRead : 1'b0)));
  assign _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowWrite = (((_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute ? execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_allowWrite : 1'b0) | (_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_1 ? execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_allowWrite : 1'b0)) | ((_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_2 ? execute_ctrl3_down_MMU_L0_ENTRIES_lane0_2_allowWrite : 1'b0) | (_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_3 ? execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_allowWrite : 1'b0)));
  assign _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowUser = (((_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute ? execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_allowUser : 1'b0) | (_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_1 ? execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_allowUser : 1'b0)) | ((_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_2 ? execute_ctrl3_down_MMU_L0_ENTRIES_lane0_2_allowUser : 1'b0) | (_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_3 ? execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_allowUser : 1'b0)));
  assign _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_3 = (((_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute ? fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_allowExecute : 1'b0) | (_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_1 ? fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_allowExecute : 1'b0)) | (_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_2 ? fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_allowExecute : 1'b0));
  assign _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowRead = (((_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute ? fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_allowRead : 1'b0) | (_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_1 ? fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_allowRead : 1'b0)) | (_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_2 ? fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_allowRead : 1'b0));
  assign _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowWrite = (((_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute ? fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_allowWrite : 1'b0) | (_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_1 ? fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_allowWrite : 1'b0)) | (_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_2 ? fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_allowWrite : 1'b0));
  assign _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowUser = (((_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute ? fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_allowUser : 1'b0) | (_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_1 ? fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_allowUser : 1'b0)) | (_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_2 ? fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_allowUser : 1'b0));
  assign _zz_MmuPlugin_logic_refill_load_nextLevelBase = MmuPlugin_logic_refill_load_readed[53 : 28];
  assign _zz_bits_pte_ppn = MmuPlugin_logic_refill_load_readed[63 : 10];
  assign _zz_PerformanceCounterPlugin_logic_fsm_calc_a = PerformanceCounterPlugin_logic_fsm_counterReaded[6:0];
  assign _zz_PerformanceCounterPlugin_logic_fsm_calc_sum_1 = {1'b0,PerformanceCounterPlugin_logic_fsm_calc_b};
  assign _zz_PerformanceCounterPlugin_logic_fsm_calc_sum = {56'd0, _zz_PerformanceCounterPlugin_logic_fsm_calc_sum_1};
  assign _zz_PerformanceCounterPlugin_logic_flusher_hits_ohFirst_masked = (PerformanceCounterPlugin_logic_flusher_hits_ohFirst_input - 2'b01);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_35 = ({19'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue ? MmuPlugin_logic_status_mxr : 1'b0)} <<< 5'd19);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_34 = {44'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_35};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_37 = ({18'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue ? MmuPlugin_logic_status_sum : 1'b0)} <<< 5'd18);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_36 = {45'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_37};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_40 = ({19'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_1 ? MmuPlugin_logic_status_mxr : 1'b0)} <<< 5'd19);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_39 = {44'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_40};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_42 = ({18'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_1 ? MmuPlugin_logic_status_sum : 1'b0)} <<< 5'd18);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_41 = {45'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_42};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_45 = ({60'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_2 ? MmuPlugin_logic_satp_mode : 4'b0000)} <<< 6'd60);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_47 = 44'h0;
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_46 = {20'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_47};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_50 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_2 ? MmuPlugin_logic_satp_ppn : 44'h0);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_49 = {20'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_50};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_52 = ({10'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3 ? PmpPlugin_logic_entries_0_address[20 : 1] : 20'h0)} <<< 4'd10);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_51 = {34'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_52};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_56 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3 ? _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4 : 10'h0);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_55 = {54'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_56};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_58 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5 ? PmpPlugin_logic_entries_0_cfg_read : 1'b0);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_57 = {63'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_58};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_61 = ({1'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5 ? PmpPlugin_logic_entries_0_cfg_write : 1'b0)} <<< 1'd1);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_60 = {62'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_61};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_63 = ({2'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5 ? PmpPlugin_logic_entries_0_cfg_execute : 1'b0)} <<< 2'd2);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_62 = {61'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_63};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_67 = ({3'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5 ? PmpPlugin_logic_entries_0_cfg_kind : 2'b00)} <<< 2'd3);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_66 = {59'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_67};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_69 = ({7'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5 ? PmpPlugin_logic_entries_0_cfg_locked : 1'b0)} <<< 3'd7);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_68 = {56'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_69};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_72 = ({10'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_6 ? PmpPlugin_logic_entries_1_address[20 : 1] : 20'h0)} <<< 4'd10);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_71 = {34'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_72};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_74 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_6 ? _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_7 : 10'h0);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_73 = {54'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_74};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_78 = ({8'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5 ? PmpPlugin_logic_entries_1_cfg_read : 1'b0)} <<< 4'd8);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_77 = {55'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_78};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_80 = ({9'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5 ? PmpPlugin_logic_entries_1_cfg_write : 1'b0)} <<< 4'd9);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_79 = {54'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_80};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_83 = ({10'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5 ? PmpPlugin_logic_entries_1_cfg_execute : 1'b0)} <<< 4'd10);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_82 = {53'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_83};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_85 = ({11'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5 ? PmpPlugin_logic_entries_1_cfg_kind : 2'b00)} <<< 4'd11);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_84 = {51'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_85};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_89 = ({15'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5 ? PmpPlugin_logic_entries_1_cfg_locked : 1'b0)} <<< 4'd15);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_88 = {48'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_89};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_91 = ({10'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_8 ? PmpPlugin_logic_entries_2_address[20 : 1] : 20'h0)} <<< 4'd10);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_90 = {34'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_91};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_94 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_8 ? _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_9 : 10'h0);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_93 = {54'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_94};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_96 = ({16'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5 ? PmpPlugin_logic_entries_2_cfg_read : 1'b0)} <<< 5'd16);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_95 = {47'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_96};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_100 = ({17'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5 ? PmpPlugin_logic_entries_2_cfg_write : 1'b0)} <<< 5'd17);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_99 = {46'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_100};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_102 = ({18'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5 ? PmpPlugin_logic_entries_2_cfg_execute : 1'b0)} <<< 5'd18);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_101 = {45'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_102};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_105 = ({19'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5 ? PmpPlugin_logic_entries_2_cfg_kind : 2'b00)} <<< 5'd19);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_104 = {43'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_105};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_107 = ({23'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5 ? PmpPlugin_logic_entries_2_cfg_locked : 1'b0)} <<< 5'd23);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_106 = {40'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_107};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_111 = ({10'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_10 ? PmpPlugin_logic_entries_3_address[20 : 1] : 20'h0)} <<< 4'd10);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_110 = {34'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_111};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_113 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_10 ? _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_11 : 10'h0);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_112 = {54'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_113};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_116 = ({24'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5 ? PmpPlugin_logic_entries_3_cfg_read : 1'b0)} <<< 5'd24);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_115 = {39'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_116};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_118 = ({25'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5 ? PmpPlugin_logic_entries_3_cfg_write : 1'b0)} <<< 5'd25);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_117 = {38'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_118};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_122 = ({26'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5 ? PmpPlugin_logic_entries_3_cfg_execute : 1'b0)} <<< 5'd26);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_121 = {37'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_122};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_124 = ({27'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5 ? PmpPlugin_logic_entries_3_cfg_kind : 2'b00)} <<< 5'd27);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_123 = {35'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_124};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_127 = ({31'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5 ? PmpPlugin_logic_entries_3_cfg_locked : 1'b0)} <<< 5'd31);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_126 = {32'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_127};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_131 = ((when_CsrService_l232 && REG_CSR_3858) ? 6'h2e : 6'h0);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_130 = {58'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_131};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_136 = ({7'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_12 ? PrivilegedPlugin_logic_harts_0_m_status_mpie : 1'b0)} <<< 3'd7);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_135 = {56'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_136};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_138 = ({3'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_12 ? PrivilegedPlugin_logic_harts_0_m_status_mie : 1'b0)} <<< 2'd3);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_137 = {60'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_138};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_141 = ({11'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_12 ? PrivilegedPlugin_logic_harts_0_m_status_mpp : 2'b00)} <<< 4'd11);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_140 = {51'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_141};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_142 = ({63'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_12 ? PrivilegedPlugin_logic_harts_0_m_status_sd : 1'b0)} <<< 6'd63);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_146 = ({17'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_12 ? PrivilegedPlugin_logic_harts_0_m_status_mprv : 1'b0)} <<< 5'd17);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_145 = {46'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_146};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_148 = ({13'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_12 ? PrivilegedPlugin_logic_harts_0_m_status_fs : 2'b00)} <<< 4'd13);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_147 = {49'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_148};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_151 = ({32'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_12 ? 2'b10 : 2'b00)} <<< 6'd32);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_150 = {30'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_151};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_153 = ({34'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_12 ? 2'b10 : 2'b00)} <<< 6'd34);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_152 = {28'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_153};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_157 = ({22'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_12 ? PrivilegedPlugin_logic_harts_0_m_status_tsr : 1'b0)} <<< 5'd22);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_156 = {41'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_157};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_159 = ({20'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_12 ? PrivilegedPlugin_logic_harts_0_m_status_tvm : 1'b0)} <<< 5'd20);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_158 = {43'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_159};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_162 = ({21'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_12 ? PrivilegedPlugin_logic_harts_0_m_status_tw : 1'b0)} <<< 5'd21);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_161 = {42'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_162};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_163 = ({63'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_13 ? PrivilegedPlugin_logic_harts_0_m_cause_interrupt : 1'b0)} <<< 6'd63);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_167 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_13 ? PrivilegedPlugin_logic_harts_0_m_cause_code : 4'b0000);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_166 = {60'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_167};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_169 = ({11'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_15 ? PrivilegedPlugin_logic_harts_0_m_ip_meip : 1'b0)} <<< 4'd11);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_168 = {52'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_169};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_172 = ({7'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_15 ? PrivilegedPlugin_logic_harts_0_m_ip_mtip : 1'b0)} <<< 3'd7);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_171 = {56'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_172};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_174 = ({3'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_15 ? PrivilegedPlugin_logic_harts_0_m_ip_msip : 1'b0)} <<< 2'd3);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_173 = {60'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_174};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_178 = ({11'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_17 ? PrivilegedPlugin_logic_harts_0_m_ie_meie : 1'b0)} <<< 4'd11);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_177 = {52'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_178};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_180 = ({7'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_17 ? PrivilegedPlugin_logic_harts_0_m_ie_mtie : 1'b0)} <<< 3'd7);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_179 = {56'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_180};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_183 = ({3'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_17 ? PrivilegedPlugin_logic_harts_0_m_ie_msie : 1'b0)} <<< 2'd3);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_182 = {60'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_183};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_185 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_18 ? PrivilegedPlugin_logic_harts_0_m_edeleg_iam : 1'b0);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_184 = {63'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_185};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_189 = ({3'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_18 ? PrivilegedPlugin_logic_harts_0_m_edeleg_bp : 1'b0)} <<< 2'd3);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_188 = {60'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_189};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_191 = ({8'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_18 ? PrivilegedPlugin_logic_harts_0_m_edeleg_eu : 1'b0)} <<< 4'd8);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_190 = {55'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_191};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_194 = ({9'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_18 ? PrivilegedPlugin_logic_harts_0_m_edeleg_es : 1'b0)} <<< 4'd9);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_193 = {54'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_194};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_196 = ({12'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_18 ? PrivilegedPlugin_logic_harts_0_m_edeleg_ipf : 1'b0)} <<< 4'd12);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_195 = {51'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_196};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_200 = ({13'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_18 ? PrivilegedPlugin_logic_harts_0_m_edeleg_lpf : 1'b0)} <<< 4'd13);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_199 = {50'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_200};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_202 = ({15'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_18 ? PrivilegedPlugin_logic_harts_0_m_edeleg_spf : 1'b0)} <<< 4'd15);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_201 = {48'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_202};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_205 = ({9'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_20 ? PrivilegedPlugin_logic_harts_0_m_ideleg_se : 1'b0)} <<< 4'd9);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_204 = {54'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_205};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_207 = ({5'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_20 ? PrivilegedPlugin_logic_harts_0_m_ideleg_st : 1'b0)} <<< 3'd5);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_206 = {58'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_207};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_211 = ({1'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_20 ? PrivilegedPlugin_logic_harts_0_m_ideleg_ss : 1'b0)} <<< 1'd1);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_210 = {62'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_211};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_213 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_21 ? PrivilegedPlugin_logic_harts_0_m_topi_priority : 1'b0);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_212 = {63'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_213};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_216 = ({16'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_21 ? PrivilegedPlugin_logic_harts_0_m_topi_interrupt : 4'b0000)} <<< 5'd16);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_215 = {44'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_216};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_218 = ({1'd0,((when_CsrService_l232 && _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_22) ? PrivilegedPlugin_logic_harts_0_mcounteren_tm : 1'b0)} <<< 1'd1);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_217 = {62'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_218};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_221 = ({63'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_23 ? PrivilegedPlugin_logic_harts_0_s_cause_interrupt : 1'b0)} <<< 6'd63);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_223 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_23 ? PrivilegedPlugin_logic_harts_0_s_cause_code : 4'b0000);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_222 = {60'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_223};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_225 = ({63'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_24 ? PrivilegedPlugin_logic_harts_0_m_status_sd : 1'b0)} <<< 6'd63);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_227 = ({8'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_12 ? PrivilegedPlugin_logic_harts_0_s_status_spp : 1'b0)} <<< 4'd8);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_226 = {55'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_227};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_231 = ({5'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_12 ? PrivilegedPlugin_logic_harts_0_s_status_spie : 1'b0)} <<< 3'd5);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_230 = {58'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_231};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_233 = ({1'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_12 ? PrivilegedPlugin_logic_harts_0_s_status_sie : 1'b0)} <<< 1'd1);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_232 = {62'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_233};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_236 = ({8'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_24 ? PrivilegedPlugin_logic_harts_0_s_status_spp : 1'b0)} <<< 4'd8);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_235 = {55'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_236};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_238 = ({5'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_24 ? PrivilegedPlugin_logic_harts_0_s_status_spie : 1'b0)} <<< 3'd5);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_237 = {58'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_238};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_242 = ({1'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_24 ? PrivilegedPlugin_logic_harts_0_s_status_sie : 1'b0)} <<< 1'd1);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_241 = {62'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_242};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_244 = ({32'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_24 ? 2'b10 : 2'b00)} <<< 6'd32);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_243 = {30'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_244};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_246 = ({63'd0,((when_CsrService_l232 && _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_25) ? PrivilegedPlugin_logic_harts_0_s_sstc_envcfg_enable : 1'b0)} <<< 6'd63);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_248 = ({13'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_24 ? PrivilegedPlugin_logic_harts_0_m_status_fs : 2'b00)} <<< 4'd13);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_247 = {49'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_248};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_252 = ({9'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_26 ? (PrivilegedPlugin_logic_harts_0_s_ie_seie && PrivilegedPlugin_logic_harts_0_m_ideleg_se) : 1'b0)} <<< 4'd9);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_251 = {54'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_252};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_254 = ({5'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_26 ? (PrivilegedPlugin_logic_harts_0_s_ie_stie && PrivilegedPlugin_logic_harts_0_m_ideleg_st) : 1'b0)} <<< 3'd5);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_253 = {58'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_254};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_257 = ({1'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_26 ? (PrivilegedPlugin_logic_harts_0_s_ie_ssie && PrivilegedPlugin_logic_harts_0_m_ideleg_ss) : 1'b0)} <<< 1'd1);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_256 = {62'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_257};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_259 = ({9'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_27 ? (PrivilegedPlugin_logic_harts_0_s_ip_seipOr && PrivilegedPlugin_logic_harts_0_m_ideleg_se) : 1'b0)} <<< 4'd9);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_258 = {54'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_259};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_263 = ({1'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_27 ? (PrivilegedPlugin_logic_harts_0_s_ip_ssip && PrivilegedPlugin_logic_harts_0_m_ideleg_ss) : 1'b0)} <<< 1'd1);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_262 = {62'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_263};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_265 = ({9'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_17 ? PrivilegedPlugin_logic_harts_0_s_ie_seie : 1'b0)} <<< 4'd9);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_264 = {54'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_265};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_268 = ({5'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_17 ? PrivilegedPlugin_logic_harts_0_s_ie_stie : 1'b0)} <<< 3'd5);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_267 = {58'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_268};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_270 = ({1'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_17 ? PrivilegedPlugin_logic_harts_0_s_ie_ssie : 1'b0)} <<< 1'd1);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_269 = {62'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_270};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_274 = ({9'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_15 ? PrivilegedPlugin_logic_harts_0_s_ip_seipOr : 1'b0)} <<< 4'd9);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_273 = {54'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_274};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_276 = ({5'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_15 ? PrivilegedPlugin_logic_harts_0_s_ip_stipOr : 1'b0)} <<< 3'd5);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_275 = {58'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_276};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_279 = ({5'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_27 ? (PrivilegedPlugin_logic_harts_0_s_ip_stipOr && PrivilegedPlugin_logic_harts_0_m_ideleg_st) : 1'b0)} <<< 3'd5);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_278 = {58'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_279};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_281 = ({1'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_15 ? PrivilegedPlugin_logic_harts_0_s_ip_ssip : 1'b0)} <<< 1'd1);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_280 = {62'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_281};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_285 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_28 ? PrivilegedPlugin_logic_harts_0_s_topi_priority : 1'b0);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_284 = {63'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_285};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_287 = ({16'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_28 ? PrivilegedPlugin_logic_harts_0_s_topi_interrupt : 4'b0000)} <<< 5'd16);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_286 = {44'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_287};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_290 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_22 ? PerformanceCounterPlugin_logic_counters_cycle_mcounteren : 1'b0);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_289 = {63'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_290};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_294 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_29 ? PerformanceCounterPlugin_logic_counters_cycle_scounteren : 1'b0);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_293 = {63'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_294};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_296 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_30 ? PerformanceCounterPlugin_logic_counters_cycle_mcountinhibit : 1'b0);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_295 = {63'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_296};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_299 = ({2'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_22 ? PerformanceCounterPlugin_logic_counters_instret_mcounteren : 1'b0)} <<< 2'd2);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_298 = {61'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_299};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_301 = ({2'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_29 ? PerformanceCounterPlugin_logic_counters_instret_scounteren : 1'b0)} <<< 2'd2);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_300 = {61'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_301};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_305 = ({2'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_30 ? PerformanceCounterPlugin_logic_counters_instret_mcountinhibit : 1'b0)} <<< 2'd2);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_304 = {61'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_305};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_307 = ({4'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_25 ? LsuPlugin_logic_cbmCsr_menvcfg_cbie : 2'b00)} <<< 3'd4);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_306 = {58'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_307};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_310 = ({6'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_25 ? LsuPlugin_logic_cbmCsr_menvcfg_cbcfe : 1'b0)} <<< 3'd6);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_309 = {57'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_310};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_312 = ({4'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_31 ? LsuPlugin_logic_cbmCsr_senvcfg_cbie : 2'b00)} <<< 3'd4);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_311 = {58'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_312};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_316 = ({6'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_31 ? LsuPlugin_logic_cbmCsr_senvcfg_cbcfe : 1'b0)} <<< 3'd6);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_315 = {57'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_316};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_319 = ({13'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_14 ? PerformanceCounterPlugin_logic_interrupt_ip : 1'b0)} <<< 4'd13);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_318 = {50'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_319};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_321 = ({13'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_16 ? PerformanceCounterPlugin_logic_interrupt_ie : 1'b0)} <<< 4'd13);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_320 = {50'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_321};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_323 = ({13'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_19 ? PerformanceCounterPlugin_logic_interrupt_sup_deleg : 1'b0)} <<< 4'd13);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_322 = {50'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_323};
  assign _zz_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask_1 = CsrAccessPlugin_logic_fsm_interface_uop[19 : 15];
  assign _zz_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask = {59'd0, _zz_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask_1};
  assign _zz_CsrRamPlugin_logic_writeLogic_hits_ohFirst_masked = (CsrRamPlugin_logic_writeLogic_hits_ohFirst_input - 4'b0001);
  assign _zz_CsrRamPlugin_logic_readLogic_hits_ohFirst_masked = (CsrRamPlugin_logic_readLogic_hits_ohFirst_input - 3'b001);
  assign _zz_CsrRamPlugin_logic_flush_counter_1 = (! CsrRamPlugin_logic_flush_done);
  assign _zz_CsrRamPlugin_logic_flush_counter = {4'd0, _zz_CsrRamPlugin_logic_flush_counter_1};
  assign _zz_execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0_1 = _zz_execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0_2[0];
  assign _zz_execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0_2 = (|{((execute_lane0_logic_decoding_decodingBits & 32'h00002030) == 32'h00002010),{_zz_execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0,{((execute_lane0_logic_decoding_decodingBits & 32'h00001030) == 32'h00000010),{((execute_lane0_logic_decoding_decodingBits & 32'h02002050) == 32'h00002010),((execute_lane0_logic_decoding_decodingBits & 32'h02001050) == 32'h00000010)}}}});
  assign _zz_execute_ctrl1_down_early0_BarrelShifterPlugin_SEL_lane0 = _zz_execute_ctrl1_down_early0_BarrelShifterPlugin_SEL_lane0_1[0];
  assign _zz_execute_ctrl1_down_early0_BarrelShifterPlugin_SEL_lane0_1 = (|{((execute_lane0_logic_decoding_decodingBits & 32'h00003034) == 32'h00001010),((execute_lane0_logic_decoding_decodingBits & 32'h02003054) == 32'h00001010)});
  assign _zz_execute_ctrl1_down_early0_BranchPlugin_SEL_lane0 = _zz_execute_ctrl1_down_early0_BranchPlugin_SEL_lane0_1[0];
  assign _zz_execute_ctrl1_down_early0_BranchPlugin_SEL_lane0_1 = (|_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0);
  assign _zz_execute_ctrl1_down_early0_MulPlugin_SEL_lane0 = _zz_execute_ctrl1_down_early0_MulPlugin_SEL_lane0_1[0];
  assign _zz_execute_ctrl1_down_early0_MulPlugin_SEL_lane0_1 = (|((execute_lane0_logic_decoding_decodingBits & 32'h02004074) == 32'h02000030));
  assign _zz_execute_ctrl1_down_early0_DivPlugin_SEL_lane0 = _zz_execute_ctrl1_down_early0_DivPlugin_SEL_lane0_1[0];
  assign _zz_execute_ctrl1_down_early0_DivPlugin_SEL_lane0_1 = (|_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0);
  assign _zz_execute_ctrl1_down_early0_EnvPlugin_SEL_lane0 = _zz_execute_ctrl1_down_early0_EnvPlugin_SEL_lane0_1[0];
  assign _zz_execute_ctrl1_down_early0_EnvPlugin_SEL_lane0_1 = (|{((execute_lane0_logic_decoding_decodingBits & 32'h00003050) == 32'h00000050),((execute_lane0_logic_decoding_decodingBits & 32'h00003058) == 32'h00001008)});
  assign _zz_execute_ctrl1_down_MulPlugin_HIGH_lane0 = _zz_execute_ctrl1_down_MulPlugin_HIGH_lane0_1[0];
  assign _zz_execute_ctrl1_down_MulPlugin_HIGH_lane0_1 = (|{((execute_lane0_logic_decoding_decodingBits & 32'h02006074) == 32'h02002030),((execute_lane0_logic_decoding_decodingBits & 32'h02005074) == 32'h02001030)});
  assign _zz_execute_ctrl1_down_CsrAccessPlugin_SEL_lane0 = _zz_execute_ctrl1_down_CsrAccessPlugin_SEL_lane0_1[0];
  assign _zz_execute_ctrl1_down_CsrAccessPlugin_SEL_lane0_1 = (|{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0_2,_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0_1});
  assign _zz_execute_ctrl1_down_AguPlugin_SEL_lane0 = _zz_execute_ctrl1_down_AguPlugin_SEL_lane0_1[0];
  assign _zz_execute_ctrl1_down_AguPlugin_SEL_lane0_1 = (|{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_2,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_1,_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0}});
  assign _zz_execute_ctrl1_down_LsuPlugin_logic_FENCE_lane0 = _zz_execute_ctrl1_down_LsuPlugin_logic_FENCE_lane0_1[0];
  assign _zz_execute_ctrl1_down_LsuPlugin_logic_FENCE_lane0_1 = (|((execute_lane0_logic_decoding_decodingBits & 32'h00003058) == 32'h00000008));
  assign _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0 = _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_1[0];
  assign _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_1 = (|{_zz_execute_ctrl1_down_AguPlugin_ATOMIC_lane0,{((execute_lane0_logic_decoding_decodingBits & 32'h00001010) == 32'h00001010),{((execute_lane0_logic_decoding_decodingBits & 32'h00002010) == 32'h00002010),{((execute_lane0_logic_decoding_decodingBits & 32'h00000050) == 32'h00000010),{_zz_execute_ctrl1_down_BYPASSED_AT_3_lane0,_zz_execute_ctrl1_down_AguPlugin_LOAD_lane0}}}}});
  assign _zz_execute_ctrl1_down_COMPLETION_AT_2_lane0 = _zz_execute_ctrl1_down_COMPLETION_AT_2_lane0_1[0];
  assign _zz_execute_ctrl1_down_COMPLETION_AT_2_lane0_1 = (|{_zz_execute_ctrl1_down_BYPASSED_AT_3_lane0_1,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0,{_zz_execute_ctrl1_down_BYPASSED_AT_3_lane0,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_3,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_2,_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_1}}}}});
  assign _zz_execute_ctrl1_down_COMPLETION_AT_4_lane0 = _zz_execute_ctrl1_down_COMPLETION_AT_4_lane0_1[0];
  assign _zz_execute_ctrl1_down_COMPLETION_AT_4_lane0_1 = (|{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_2,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_1,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0,_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_3}}});
  assign _zz_execute_ctrl1_down_COMPLETION_AT_3_lane0 = _zz_execute_ctrl1_down_COMPLETION_AT_3_lane0_1[0];
  assign _zz_execute_ctrl1_down_COMPLETION_AT_3_lane0_1 = (|{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0_2,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0_1,_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0}});
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_4 = _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_5[0];
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_5 = (|{_zz_execute_ctrl1_down_BYPASSED_AT_3_lane0_1,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0,{_zz_execute_ctrl1_down_BYPASSED_AT_3_lane0,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_3,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_2,_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_1}}}}});
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_4 = _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_5[0];
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_5 = (|{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_2,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_1,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0,_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_3}}});
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0_3 = _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0_4[0];
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0_4 = (|{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0_2,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0_1,_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0}});
  assign _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0_1 = _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0_2[0];
  assign _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0_2 = (|{_zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0,_zz_execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0});
  assign _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_SLTX_lane0 = _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_SLTX_lane0_1[0];
  assign _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_SLTX_lane0_1 = (|((execute_lane0_logic_decoding_decodingBits & 32'h00006004) == 32'h00002000));
  assign _zz_execute_ctrl1_down_SrcStageables_REVERT_lane0 = _zz_execute_ctrl1_down_SrcStageables_REVERT_lane0_1[0];
  assign _zz_execute_ctrl1_down_SrcStageables_REVERT_lane0_1 = (|{_zz_execute_ctrl1_down_BYPASSED_AT_3_lane0_2,{((execute_lane0_logic_decoding_decodingBits & 32'h00002014) == 32'h00002010),((execute_lane0_logic_decoding_decodingBits & 32'h40000034) == 32'h40000030)}});
  assign _zz_execute_ctrl1_down_SrcStageables_ZERO_lane0 = _zz_execute_ctrl1_down_SrcStageables_ZERO_lane0_1[0];
  assign _zz_execute_ctrl1_down_SrcStageables_ZERO_lane0_1 = (|{((execute_lane0_logic_decoding_decodingBits & 32'h00000024) == 32'h00000024),((execute_lane0_logic_decoding_decodingBits & 32'h00000018) == 32'h00000008)});
  assign _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_SIGNED_lane0 = _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_SIGNED_lane0_1[0];
  assign _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_SIGNED_lane0_1 = (|{_zz_execute_ctrl1_down_RsUnsignedPlugin_IS_W_lane0,((execute_lane0_logic_decoding_decodingBits & 32'h00004010) == 32'h0)});
  assign _zz_execute_ctrl1_down_BYPASSED_AT_2_lane0 = _zz_execute_ctrl1_down_BYPASSED_AT_2_lane0_1[0];
  assign _zz_execute_ctrl1_down_BYPASSED_AT_2_lane0_1 = (|{_zz_execute_ctrl1_down_BYPASSED_AT_3_lane0_1,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0,{_zz_execute_ctrl1_down_BYPASSED_AT_3_lane0,{((execute_lane0_logic_decoding_decodingBits & 32'h02000068) == 32'h00000020),((execute_lane0_logic_decoding_decodingBits & 32'h02002060) == 32'h00000020)}}}});
  assign _zz_execute_ctrl1_down_BYPASSED_AT_3_lane0_3 = _zz_execute_ctrl1_down_BYPASSED_AT_3_lane0_4[0];
  assign _zz_execute_ctrl1_down_BYPASSED_AT_3_lane0_4 = (|{_zz_execute_ctrl1_down_BYPASSED_AT_3_lane0_2,{((execute_lane0_logic_decoding_decodingBits & 32'h00004020) == 32'h00004020),{_zz_execute_ctrl1_down_BYPASSED_AT_3_lane0_1,{_zz_execute_ctrl1_down_BYPASSED_AT_3_lane0,{((execute_lane0_logic_decoding_decodingBits & 32'h02002020) == 32'h00000020),((execute_lane0_logic_decoding_decodingBits & 32'h02000028) == 32'h00000020)}}}}});
  assign _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane0 = _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane0_1[0];
  assign _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane0_1 = (|{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_2,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_1,_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0}});
  assign _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane0 = _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane0_1[0];
  assign _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane0_1 = (|{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_2,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_1,_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0}});
  assign _zz_execute_ctrl1_down_SrcStageables_UNSIGNED_lane0 = _zz_execute_ctrl1_down_SrcStageables_UNSIGNED_lane0_1[0];
  assign _zz_execute_ctrl1_down_SrcStageables_UNSIGNED_lane0_1 = (|{((execute_lane0_logic_decoding_decodingBits & 32'h00002010) == 32'h00002000),((execute_lane0_logic_decoding_decodingBits & 32'h00005000) == 32'h00001000)});
  assign _zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0_1 = _zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0_2[0];
  assign _zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0_2 = (|_zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0);
  assign _zz_execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane0 = _zz_execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane0_1[0];
  assign _zz_execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane0_1 = (|((execute_lane0_logic_decoding_decodingBits & 32'h40000000) == 32'h40000000));
  assign _zz_execute_ctrl1_down_BarrelShifterPlugin_IS_W_lane0 = _zz_execute_ctrl1_down_BarrelShifterPlugin_IS_W_lane0_1[0];
  assign _zz_execute_ctrl1_down_BarrelShifterPlugin_IS_W_lane0_1 = (|_zz_execute_ctrl1_down_RsUnsignedPlugin_IS_W_lane0);
  assign _zz_execute_ctrl1_down_BarrelShifterPlugin_IS_W_RIGHT_lane0 = _zz_execute_ctrl1_down_BarrelShifterPlugin_IS_W_RIGHT_lane0_1[0];
  assign _zz_execute_ctrl1_down_BarrelShifterPlugin_IS_W_RIGHT_lane0_1 = (|((execute_lane0_logic_decoding_decodingBits & 32'h00004008) == 32'h00004008));
  assign _zz_execute_ctrl1_down_RsUnsignedPlugin_RS1_SIGNED_lane0 = _zz_execute_ctrl1_down_RsUnsignedPlugin_RS1_SIGNED_lane0_1[0];
  assign _zz_execute_ctrl1_down_RsUnsignedPlugin_RS1_SIGNED_lane0_1 = (|{((execute_lane0_logic_decoding_decodingBits & 32'h00001000) == 32'h0),_zz_execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0});
  assign _zz_execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0_1 = _zz_execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0_2[0];
  assign _zz_execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0_2 = (|{((execute_lane0_logic_decoding_decodingBits & 32'h00005000) == 32'h00004000),_zz_execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0});
  assign _zz_execute_ctrl1_down_DivPlugin_REM_lane0 = _zz_execute_ctrl1_down_DivPlugin_REM_lane0_1[0];
  assign _zz_execute_ctrl1_down_DivPlugin_REM_lane0_1 = (|_zz_execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0);
  assign _zz_execute_ctrl1_down_RsUnsignedPlugin_IS_W_lane0_1 = _zz_execute_ctrl1_down_RsUnsignedPlugin_IS_W_lane0_2[0];
  assign _zz_execute_ctrl1_down_RsUnsignedPlugin_IS_W_lane0_2 = (|_zz_execute_ctrl1_down_RsUnsignedPlugin_IS_W_lane0);
  assign _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_IMM_lane0 = _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_IMM_lane0_1[0];
  assign _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_IMM_lane0_1 = (|((execute_lane0_logic_decoding_decodingBits & 32'h00004000) == 32'h00004000));
  assign _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0_1 = _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0_2[0];
  assign _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0_2 = (|_zz_execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0);
  assign _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0_1 = _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0_2[0];
  assign _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0_2 = (|_zz_execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0);
  assign _zz_execute_ctrl1_down_AguPlugin_LOAD_lane0_1 = _zz_execute_ctrl1_down_AguPlugin_LOAD_lane0_2[0];
  assign _zz_execute_ctrl1_down_AguPlugin_LOAD_lane0_2 = (|{_zz_execute_ctrl1_down_AguPlugin_LOAD_lane0,{((execute_lane0_logic_decoding_decodingBits & 32'h10000028) == 32'h00000028),((execute_lane0_logic_decoding_decodingBits & 32'h18002008) == 32'h10002008)}});
  assign _zz_execute_ctrl1_down_AguPlugin_STORE_lane0_1 = _zz_execute_ctrl1_down_AguPlugin_STORE_lane0_2[0];
  assign _zz_execute_ctrl1_down_AguPlugin_STORE_lane0_2 = (|{((execute_lane0_logic_decoding_decodingBits & 32'h08000020) == 32'h08000020),{_zz_execute_ctrl1_down_AguPlugin_STORE_lane0,((execute_lane0_logic_decoding_decodingBits & 32'h00000028) == 32'h00000020)}});
  assign _zz_execute_ctrl1_down_AguPlugin_ATOMIC_lane0_1 = _zz_execute_ctrl1_down_AguPlugin_ATOMIC_lane0_2[0];
  assign _zz_execute_ctrl1_down_AguPlugin_ATOMIC_lane0_2 = (|_zz_execute_ctrl1_down_AguPlugin_ATOMIC_lane0);
  assign _zz_execute_ctrl1_down_AguPlugin_FLOAT_lane0 = _zz_execute_ctrl1_down_AguPlugin_FLOAT_lane0_1[0];
  assign _zz_execute_ctrl1_down_AguPlugin_FLOAT_lane0_1 = 1'b0;
  assign _zz_execute_ctrl1_down_AguPlugin_CLEAN_lane0 = _zz_execute_ctrl1_down_AguPlugin_CLEAN_lane0_1[0];
  assign _zz_execute_ctrl1_down_AguPlugin_CLEAN_lane0_1 = (|{((execute_lane0_logic_decoding_decodingBits & 32'h00102028) == 32'h00102008),((execute_lane0_logic_decoding_decodingBits & 32'h00202028) == 32'h00202008)});
  assign _zz_execute_ctrl1_down_AguPlugin_INVALIDATE_lane0 = _zz_execute_ctrl1_down_AguPlugin_INVALIDATE_lane0_1[0];
  assign _zz_execute_ctrl1_down_AguPlugin_INVALIDATE_lane0_1 = (|((execute_lane0_logic_decoding_decodingBits & 32'h00102028) == 32'h00002008));
  assign _zz_execute_ctrl1_down_LsuPlugin_logic_LSU_PREFETCH_lane0 = _zz_execute_ctrl1_down_LsuPlugin_logic_LSU_PREFETCH_lane0_1[0];
  assign _zz_execute_ctrl1_down_LsuPlugin_logic_LSU_PREFETCH_lane0_1 = 1'b0;
  assign _zz_WhiteboxerPlugin_logic_csr_access_payload_address = CsrAccessPlugin_logic_fsm_interface_uop;
  assign _zz__zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_1_1 = _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter;
  assign _zz__zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_1 = {59'd0, _zz__zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_1_1};
  assign _zz__zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_1_1 = _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter;
  assign _zz__zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_1 = {59'd0, _zz__zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_1_1};
  assign _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_1_1 = _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0;
  assign _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_1 = {59'd0, _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_1_1};
  assign _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_1_1 = _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1;
  assign _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_1 = {59'd0, _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_1_1};
  assign _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_1_1 = _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0;
  assign _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_1 = {59'd0, _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_1_1};
  assign _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_1_1 = _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1;
  assign _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_1 = {59'd0, _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_1_1};
  assign _zz_TrapPlugin_logic_harts_0_crsPorts_write_data_1 = TrapPlugin_logic_harts_0_trap_pending_pc;
  assign _zz_TrapPlugin_logic_harts_0_crsPorts_write_data = {{25{_zz_TrapPlugin_logic_harts_0_crsPorts_write_data_1[38]}}, _zz_TrapPlugin_logic_harts_0_crsPorts_write_data_1};
  assign _zz_TrapPlugin_logic_harts_0_crsPorts_write_data_3 = TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_tval;
  assign _zz_TrapPlugin_logic_harts_0_crsPorts_write_data_2 = {{25{_zz_TrapPlugin_logic_harts_0_crsPorts_write_data_3[38]}}, _zz_TrapPlugin_logic_harts_0_crsPorts_write_data_3};
  assign _zz_TrapPlugin_logic_harts_0_crsPorts_write_data_5 = TrapPlugin_logic_harts_0_trap_pending_pc;
  assign _zz_TrapPlugin_logic_harts_0_crsPorts_write_data_4 = {{25{_zz_TrapPlugin_logic_harts_0_crsPorts_write_data_5[38]}}, _zz_TrapPlugin_logic_harts_0_crsPorts_write_data_5};
  assign _zz_TrapPlugin_logic_harts_0_trap_pcPort_payload_pc = TrapPlugin_logic_harts_0_trap_fsm_readed;
  assign _zz_TrapPlugin_logic_harts_0_trap_pcPort_payload_pc_1 = TrapPlugin_logic_harts_0_trap_fsm_readed;
  assign _zz_MmuPlugin_logic_refill_load_address = {{MmuPlugin_logic_satp_ppn,MmuPlugin_logic_refill_arbiter_io_output_payload_address[38 : 30]},3'b000};
  assign _zz_FetchL1Plugin_logic_translationStorage_logic_sl_0_write_mask = (2'b01 <<< FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_value);
  assign _zz_FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_physicalAddress = (MmuPlugin_logic_refill_load_levelToPhysicalAddress_0 >>> 4'd12);
  assign _zz_LsuPlugin_logic_translationStorage_logic_sl_0_write_mask = (MmuPlugin_logic_refill_storageOhReg[1] ? _zz_LsuPlugin_logic_translationStorage_logic_sl_0_write_mask_1 : 4'b0000);
  assign _zz_LsuPlugin_logic_translationStorage_logic_sl_0_write_mask_1 = (4'b0001 <<< LsuPlugin_logic_translationStorage_logic_sl_0_allocId_value);
  assign _zz_LsuPlugin_logic_translationStorage_logic_sl_0_write_data_physicalAddress = (MmuPlugin_logic_refill_load_levelToPhysicalAddress_0 >>> 4'd12);
  assign _zz_FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_physicalAddress = (MmuPlugin_logic_refill_load_levelToPhysicalAddress_1 >>> 5'd21);
  assign _zz_LsuPlugin_logic_translationStorage_logic_sl_1_write_data_physicalAddress = (MmuPlugin_logic_refill_load_levelToPhysicalAddress_1 >>> 5'd21);
  assign _zz_FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_physicalAddress_1 = (MmuPlugin_logic_refill_load_levelToPhysicalAddress_2 >>> 5'd21);
  assign _zz_LsuPlugin_logic_translationStorage_logic_sl_1_write_data_physicalAddress_1 = (MmuPlugin_logic_refill_load_levelToPhysicalAddress_2 >>> 5'd21);
  assign _zz_PerformanceCounterPlugin_logic_writePort_data = PerformanceCounterPlugin_logic_fsm_calc_sum;
  assign _zz_PerformanceCounterPlugin_logic_counters_cycle_value_2 = CsrAccessPlugin_bus_write_bits;
  assign _zz_PerformanceCounterPlugin_logic_counters_instret_value_2 = CsrAccessPlugin_bus_write_bits;
  assign _zz_BtbPlugin_logic_ras_mem_stack_port = BtbPlugin_logic_ras_write_payload_data;
  assign _zz_LsuL1Plugin_logic_ways_0_mem_port = {LsuL1Plugin_logic_waysWrite_tag_fault,{LsuL1Plugin_logic_waysWrite_tag_address,LsuL1Plugin_logic_waysWrite_tag_loaded}};
  assign _zz_LsuL1Plugin_logic_ways_0_mem_port_1 = LsuL1Plugin_logic_waysWrite_mask[0];
  assign _zz_LsuL1Plugin_logic_ways_1_mem_port = {LsuL1Plugin_logic_waysWrite_tag_fault,{LsuL1Plugin_logic_waysWrite_tag_address,LsuL1Plugin_logic_waysWrite_tag_loaded}};
  assign _zz_LsuL1Plugin_logic_ways_1_mem_port_1 = LsuL1Plugin_logic_waysWrite_mask[1];
  assign _zz_LsuL1Plugin_logic_shared_mem_port = {LsuL1Plugin_logic_shared_write_payload_data_dirty,LsuL1Plugin_logic_shared_write_payload_data_plru_0};
  assign _zz_LsuL1Plugin_logic_writeback_victimBuffer_port = LsuL1Plugin_logic_writeback_read_slotReadLast_payload_wordIndex;
  assign _zz_FetchL1Plugin_logic_ways_0_mem_port = {FetchL1Plugin_logic_waysWrite_tag_address,{FetchL1Plugin_logic_waysWrite_tag_error,FetchL1Plugin_logic_waysWrite_tag_loaded}};
  assign _zz_FetchL1Plugin_logic_ways_0_mem_port_1 = FetchL1Plugin_logic_waysWrite_mask[0];
  assign _zz_FetchL1Plugin_logic_ways_1_mem_port = {FetchL1Plugin_logic_waysWrite_tag_address,{FetchL1Plugin_logic_waysWrite_tag_error,FetchL1Plugin_logic_waysWrite_tag_loaded}};
  assign _zz_FetchL1Plugin_logic_ways_1_mem_port_1 = FetchL1Plugin_logic_waysWrite_mask[1];
  assign _zz_GSharePlugin_logic_mem_banks_0_port = {GSharePlugin_logic_mem_writes_0_payload_data_1,GSharePlugin_logic_mem_writes_0_payload_data_0};
  assign _zz_BtbPlugin_logic_mem_port = {BtbPlugin_logic_memDp_wp_payload_data_0_isPop,{BtbPlugin_logic_memDp_wp_payload_data_0_isPush,{BtbPlugin_logic_memDp_wp_payload_data_0_isBranch,{BtbPlugin_logic_memDp_wp_payload_data_0_pcTarget,{BtbPlugin_logic_memDp_wp_payload_data_0_sliceLow,BtbPlugin_logic_memDp_wp_payload_data_0_hash}}}}};
  assign _zz_FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_0_port = {FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowUser,{FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowExecute,{FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowWrite,{FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowRead,{FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_physicalAddress,{FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_virtualAddress,FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_valid}}}}}};
  assign _zz_FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_0_port_1 = FetchL1Plugin_logic_translationStorage_logic_sl_0_write_mask[0];
  assign _zz_FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_1_port = {FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowUser,{FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowExecute,{FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowWrite,{FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowRead,{FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_physicalAddress,{FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_virtualAddress,FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_valid}}}}}};
  assign _zz_FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_1_port_1 = FetchL1Plugin_logic_translationStorage_logic_sl_0_write_mask[1];
  assign _zz_FetchL1Plugin_logic_translationStorage_logic_sl_1_ways_0_port = {FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowUser,{FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowExecute,{FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowWrite,{FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowRead,{FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_physicalAddress,{FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_virtualAddress,FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_valid}}}}}};
  assign _zz_FetchL1Plugin_logic_translationStorage_logic_sl_1_ways_0_port_1 = FetchL1Plugin_logic_translationStorage_logic_sl_1_write_mask[0];
  assign _zz_LsuPlugin_logic_translationStorage_logic_sl_0_ways_0_port = {LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowUser,{LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowExecute,{LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowWrite,{LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowRead,{LsuPlugin_logic_translationStorage_logic_sl_0_write_data_physicalAddress,{LsuPlugin_logic_translationStorage_logic_sl_0_write_data_virtualAddress,LsuPlugin_logic_translationStorage_logic_sl_0_write_data_valid}}}}}};
  assign _zz_LsuPlugin_logic_translationStorage_logic_sl_0_ways_0_port_1 = LsuPlugin_logic_translationStorage_logic_sl_0_write_mask[0];
  assign _zz_LsuPlugin_logic_translationStorage_logic_sl_0_ways_1_port = {LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowUser,{LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowExecute,{LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowWrite,{LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowRead,{LsuPlugin_logic_translationStorage_logic_sl_0_write_data_physicalAddress,{LsuPlugin_logic_translationStorage_logic_sl_0_write_data_virtualAddress,LsuPlugin_logic_translationStorage_logic_sl_0_write_data_valid}}}}}};
  assign _zz_LsuPlugin_logic_translationStorage_logic_sl_0_ways_1_port_1 = LsuPlugin_logic_translationStorage_logic_sl_0_write_mask[1];
  assign _zz_LsuPlugin_logic_translationStorage_logic_sl_0_ways_2_port = {LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowUser,{LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowExecute,{LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowWrite,{LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowRead,{LsuPlugin_logic_translationStorage_logic_sl_0_write_data_physicalAddress,{LsuPlugin_logic_translationStorage_logic_sl_0_write_data_virtualAddress,LsuPlugin_logic_translationStorage_logic_sl_0_write_data_valid}}}}}};
  assign _zz_LsuPlugin_logic_translationStorage_logic_sl_0_ways_2_port_1 = LsuPlugin_logic_translationStorage_logic_sl_0_write_mask[2];
  assign _zz_LsuPlugin_logic_translationStorage_logic_sl_1_ways_0_port = {LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowUser,{LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowExecute,{LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowWrite,{LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowRead,{LsuPlugin_logic_translationStorage_logic_sl_1_write_data_physicalAddress,{LsuPlugin_logic_translationStorage_logic_sl_1_write_data_virtualAddress,LsuPlugin_logic_translationStorage_logic_sl_1_write_data_valid}}}}}};
  assign _zz_LsuPlugin_logic_translationStorage_logic_sl_1_ways_0_port_1 = LsuPlugin_logic_translationStorage_logic_sl_1_write_mask[0];
  assign _zz_57 = {_zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0_1,_zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0};
  assign _zz_59 = {_zz_22[2],{_zz_22[1],_zz_22[0]}};
  assign _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_0_1 = fetch_logic_ctrls_1_down_Fetch_WORD_PC[2 : 2];
  assign _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_1_1 = fetch_logic_ctrls_1_down_Fetch_WORD_PC[2 : 2];
  assign _zz_PerformanceCounterPlugin_logic_commitCount_1 = PerformanceCounterPlugin_logic_commitMask[0];
  assign _zz_LsuPlugin_logic_onCtrl_loadData_shifted_1 = execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0[2 : 0];
  assign _zz_LsuPlugin_logic_onCtrl_loadData_shifted_3 = execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0[2 : 1];
  assign _zz_LsuPlugin_logic_onCtrl_loadData_shifted_5 = execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0[2 : 2];
  assign _zz_LsuPlugin_logic_onCtrl_loadData_shifted_7 = execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0[2 : 2];
  assign _zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK_1 = fetch_logic_ctrls_2_down_Fetch_WORD_PC[1 : 1];
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_24 = AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 10];
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_26 = {AlignerPlugin_logic_extractors_0_ctx_instruction[12],AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 5]};
  assign _zz_PerformanceCounterPlugin_logic_events_sums_0_2 = _zz_PerformanceCounterPlugin_logic_events_sums_0[0];
  assign _zz_PerformanceCounterPlugin_logic_events_sums_1_2 = _zz_PerformanceCounterPlugin_logic_events_sums_1[0];
  assign _zz_PerformanceCounterPlugin_logic_events_sums_2_2 = _zz_PerformanceCounterPlugin_logic_events_sums_2[0];
  assign _zz_PerformanceCounterPlugin_logic_events_sums_3_2 = _zz_PerformanceCounterPlugin_logic_events_sums_3[0];
  assign _zz_PerformanceCounterPlugin_logic_events_sums_4_2 = _zz_PerformanceCounterPlugin_logic_events_sums_4[0];
  assign _zz_PerformanceCounterPlugin_logic_events_sums_5_2 = _zz_PerformanceCounterPlugin_logic_events_sums_5[0];
  assign _zz_PerformanceCounterPlugin_logic_events_sums_6_2 = _zz_PerformanceCounterPlugin_logic_events_sums_6[0];
  assign _zz_PerformanceCounterPlugin_logic_events_sums_7_2 = _zz_PerformanceCounterPlugin_logic_events_sums_7[0];
  assign _zz_PerformanceCounterPlugin_logic_events_sums_8_2 = _zz_PerformanceCounterPlugin_logic_events_sums_8[0];
  assign _zz_PerformanceCounterPlugin_logic_events_sums_9_2 = _zz_PerformanceCounterPlugin_logic_events_sums_9[0];
  assign _zz_PerformanceCounterPlugin_logic_events_sums_10_2 = _zz_PerformanceCounterPlugin_logic_events_sums_10[0];
  assign _zz_PerformanceCounterPlugin_logic_events_sums_11_2 = _zz_PerformanceCounterPlugin_logic_events_sums_11[0];
  assign _zz_PerformanceCounterPlugin_logic_events_sums_12_2 = _zz_PerformanceCounterPlugin_logic_events_sums_12[0];
  assign _zz_PerformanceCounterPlugin_logic_events_sums_13_2 = _zz_PerformanceCounterPlugin_logic_events_sums_13[0];
  assign _zz_WhiteboxerPlugin_logic_perf_candidatesCount_1 = DispatchPlugin_logic_candidates_0_ctx_valid;
  assign _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCount_1 = decode_ctrls_1_up_LANE_SEL_0;
  assign _zz_early0_BarrelShifterPlugin_logic_shift_reversed_1 = execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[9];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_reversed_2 = execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[10];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_reversed_3 = {execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[11],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[12],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[13],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[14],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[15],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[16],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[17],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[18],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[19],{_zz_early0_BarrelShifterPlugin_logic_shift_reversed_4,{_zz_early0_BarrelShifterPlugin_logic_shift_reversed_5,_zz_early0_BarrelShifterPlugin_logic_shift_reversed_6}}}}}}}}}}};
  assign _zz_early0_BarrelShifterPlugin_logic_shift_reversed_4 = execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[20];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_reversed_5 = execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[21];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_reversed_6 = {execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[22],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[23],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[24],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[25],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[26],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[27],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[28],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[29],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[30],{_zz_early0_BarrelShifterPlugin_logic_shift_reversed_7,{_zz_early0_BarrelShifterPlugin_logic_shift_reversed_8,_zz_early0_BarrelShifterPlugin_logic_shift_reversed_9}}}}}}}}}}};
  assign _zz_early0_BarrelShifterPlugin_logic_shift_reversed_7 = execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[31];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_reversed_8 = execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[32];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_reversed_9 = {execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[33],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[34],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[35],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[36],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[37],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[38],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[39],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[40],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[41],{_zz_early0_BarrelShifterPlugin_logic_shift_reversed_10,{_zz_early0_BarrelShifterPlugin_logic_shift_reversed_11,_zz_early0_BarrelShifterPlugin_logic_shift_reversed_12}}}}}}}}}}};
  assign _zz_early0_BarrelShifterPlugin_logic_shift_reversed_10 = execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[42];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_reversed_11 = execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[43];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_reversed_12 = {execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[44],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[45],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[46],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[47],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[48],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[49],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[50],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[51],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[52],{_zz_early0_BarrelShifterPlugin_logic_shift_reversed_13,{_zz_early0_BarrelShifterPlugin_logic_shift_reversed_14,_zz_early0_BarrelShifterPlugin_logic_shift_reversed_15}}}}}}}}}}};
  assign _zz_early0_BarrelShifterPlugin_logic_shift_reversed_13 = execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[53];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_reversed_14 = execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[54];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_reversed_15 = {execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[55],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[56],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[57],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[58],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[59],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[60],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[61],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[62],execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[63]}}}}}}}};
  assign _zz_early0_BarrelShifterPlugin_logic_shift_patched_1 = early0_BarrelShifterPlugin_logic_shift_shifted[9];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_patched_2 = early0_BarrelShifterPlugin_logic_shift_shifted[10];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_patched_3 = {early0_BarrelShifterPlugin_logic_shift_shifted[11],{early0_BarrelShifterPlugin_logic_shift_shifted[12],{early0_BarrelShifterPlugin_logic_shift_shifted[13],{early0_BarrelShifterPlugin_logic_shift_shifted[14],{early0_BarrelShifterPlugin_logic_shift_shifted[15],{early0_BarrelShifterPlugin_logic_shift_shifted[16],{early0_BarrelShifterPlugin_logic_shift_shifted[17],{early0_BarrelShifterPlugin_logic_shift_shifted[18],{early0_BarrelShifterPlugin_logic_shift_shifted[19],{_zz_early0_BarrelShifterPlugin_logic_shift_patched_4,{_zz_early0_BarrelShifterPlugin_logic_shift_patched_5,_zz_early0_BarrelShifterPlugin_logic_shift_patched_6}}}}}}}}}}};
  assign _zz_early0_BarrelShifterPlugin_logic_shift_patched_4 = early0_BarrelShifterPlugin_logic_shift_shifted[20];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_patched_5 = early0_BarrelShifterPlugin_logic_shift_shifted[21];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_patched_6 = {early0_BarrelShifterPlugin_logic_shift_shifted[22],{early0_BarrelShifterPlugin_logic_shift_shifted[23],{early0_BarrelShifterPlugin_logic_shift_shifted[24],{early0_BarrelShifterPlugin_logic_shift_shifted[25],{early0_BarrelShifterPlugin_logic_shift_shifted[26],{early0_BarrelShifterPlugin_logic_shift_shifted[27],{early0_BarrelShifterPlugin_logic_shift_shifted[28],{early0_BarrelShifterPlugin_logic_shift_shifted[29],{early0_BarrelShifterPlugin_logic_shift_shifted[30],{_zz_early0_BarrelShifterPlugin_logic_shift_patched_7,{_zz_early0_BarrelShifterPlugin_logic_shift_patched_8,_zz_early0_BarrelShifterPlugin_logic_shift_patched_9}}}}}}}}}}};
  assign _zz_early0_BarrelShifterPlugin_logic_shift_patched_7 = early0_BarrelShifterPlugin_logic_shift_shifted[31];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_patched_8 = early0_BarrelShifterPlugin_logic_shift_shifted[32];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_patched_9 = {early0_BarrelShifterPlugin_logic_shift_shifted[33],{early0_BarrelShifterPlugin_logic_shift_shifted[34],{early0_BarrelShifterPlugin_logic_shift_shifted[35],{early0_BarrelShifterPlugin_logic_shift_shifted[36],{early0_BarrelShifterPlugin_logic_shift_shifted[37],{early0_BarrelShifterPlugin_logic_shift_shifted[38],{early0_BarrelShifterPlugin_logic_shift_shifted[39],{early0_BarrelShifterPlugin_logic_shift_shifted[40],{early0_BarrelShifterPlugin_logic_shift_shifted[41],{_zz_early0_BarrelShifterPlugin_logic_shift_patched_10,{_zz_early0_BarrelShifterPlugin_logic_shift_patched_11,_zz_early0_BarrelShifterPlugin_logic_shift_patched_12}}}}}}}}}}};
  assign _zz_early0_BarrelShifterPlugin_logic_shift_patched_10 = early0_BarrelShifterPlugin_logic_shift_shifted[42];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_patched_11 = early0_BarrelShifterPlugin_logic_shift_shifted[43];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_patched_12 = {early0_BarrelShifterPlugin_logic_shift_shifted[44],{early0_BarrelShifterPlugin_logic_shift_shifted[45],{early0_BarrelShifterPlugin_logic_shift_shifted[46],{early0_BarrelShifterPlugin_logic_shift_shifted[47],{early0_BarrelShifterPlugin_logic_shift_shifted[48],{early0_BarrelShifterPlugin_logic_shift_shifted[49],{early0_BarrelShifterPlugin_logic_shift_shifted[50],{early0_BarrelShifterPlugin_logic_shift_shifted[51],{early0_BarrelShifterPlugin_logic_shift_shifted[52],{_zz_early0_BarrelShifterPlugin_logic_shift_patched_13,{_zz_early0_BarrelShifterPlugin_logic_shift_patched_14,_zz_early0_BarrelShifterPlugin_logic_shift_patched_15}}}}}}}}}}};
  assign _zz_early0_BarrelShifterPlugin_logic_shift_patched_13 = early0_BarrelShifterPlugin_logic_shift_shifted[53];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_patched_14 = early0_BarrelShifterPlugin_logic_shift_shifted[54];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_patched_15 = {early0_BarrelShifterPlugin_logic_shift_shifted[55],{early0_BarrelShifterPlugin_logic_shift_shifted[56],{early0_BarrelShifterPlugin_logic_shift_shifted[57],{early0_BarrelShifterPlugin_logic_shift_shifted[58],{early0_BarrelShifterPlugin_logic_shift_shifted[59],{early0_BarrelShifterPlugin_logic_shift_shifted[60],{early0_BarrelShifterPlugin_logic_shift_shifted[61],{early0_BarrelShifterPlugin_logic_shift_shifted[62],early0_BarrelShifterPlugin_logic_shift_shifted[63]}}}}}}}};
  assign _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_1 = _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH[6];
  assign _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_2 = _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH[7];
  assign _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_3 = {_zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH[8],{_zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH[9],{_zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH[10],{_zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH[11],_zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH[12]}}}};
  assign _zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0_1 = _zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0[21];
  assign _zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0_2 = (_zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0[20] != LsuPlugin_logic_onPma_addressExtension);
  assign _zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0_3 = (_zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0[19] != LsuPlugin_logic_onPma_addressExtension);
  assign _zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0_4 = {(_zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0[18] != LsuPlugin_logic_onPma_addressExtension),{(_zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0[17] != LsuPlugin_logic_onPma_addressExtension),{(_zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0[16] != LsuPlugin_logic_onPma_addressExtension),{(_zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0[15] != LsuPlugin_logic_onPma_addressExtension),{(_zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0[14] != LsuPlugin_logic_onPma_addressExtension),{(_zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0_5 != LsuPlugin_logic_onPma_addressExtension),{_zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0_6,{_zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0_7,_zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0_8}}}}}}}};
  assign _zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0_5 = _zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0[13];
  assign _zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0_6 = (_zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0[12] != LsuPlugin_logic_onPma_addressExtension);
  assign _zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0_7 = (_zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0[11] != LsuPlugin_logic_onPma_addressExtension);
  assign _zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0_8 = {(_zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0[10] != LsuPlugin_logic_onPma_addressExtension),{(_zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0[9] != LsuPlugin_logic_onPma_addressExtension),{(_zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0[8] != LsuPlugin_logic_onPma_addressExtension),{(_zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0[7] != LsuPlugin_logic_onPma_addressExtension),{(_zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0[6] != LsuPlugin_logic_onPma_addressExtension),{(_zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0_9 != LsuPlugin_logic_onPma_addressExtension),{_zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0_10,{_zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0_11,_zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0_12}}}}}}}};
  assign _zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0_9 = _zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0[5];
  assign _zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0_10 = (_zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0[4] != LsuPlugin_logic_onPma_addressExtension);
  assign _zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0_11 = (_zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0[3] != LsuPlugin_logic_onPma_addressExtension);
  assign _zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0_12 = {(_zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0[2] != LsuPlugin_logic_onPma_addressExtension),{(_zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0[1] != LsuPlugin_logic_onPma_addressExtension),(_zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0[0] != LsuPlugin_logic_onPma_addressExtension)}};
  assign _zz_execute_ctrl4_down_LsuL1_ABORD_lane0 = (! execute_ctrl4_up_LANE_SEL_lane0);
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_19 = {_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_9,AlignerPlugin_logic_extractors_0_ctx_instruction[4 : 3]};
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_20 = AlignerPlugin_logic_extractors_0_ctx_instruction[5];
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_21 = AlignerPlugin_logic_extractors_0_ctx_instruction[2];
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_27 = 7'h0;
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_28 = AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 2];
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_29 = AlignerPlugin_logic_extractors_0_ctx_instruction[12];
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_30 = AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7];
  assign _zz_LsuPlugin_logic_onPma_io_rsp_fault = 32'hf0000000;
  assign _zz_LsuPlugin_logic_onPma_io_rsp_fault_1 = (LsuPlugin_pmaBuilder_io_addressBits & 32'hf0000000);
  assign _zz_LsuPlugin_logic_onPma_io_rsp_fault_2 = 32'h10000000;
  assign _zz_LsuPlugin_logic_onPma_io_rsp_fault_3 = ((LsuPlugin_pmaBuilder_io_addressBits & 32'hf8000000) == 32'h70000000);
  assign _zz_LsuPlugin_logic_onPma_io_rsp_fault_4 = ((LsuPlugin_pmaBuilder_io_addressBits & 32'hf8000000) == 32'h80000000);
  assign _zz_LsuPlugin_logic_onPma_io_rsp_fault_5 = {((LsuPlugin_pmaBuilder_io_addressBits & 32'hf1000000) == 32'h0),{((LsuPlugin_pmaBuilder_io_addressBits & 32'hfc000000) == 32'h78000000),{((LsuPlugin_pmaBuilder_io_addressBits & 32'hfe000000) == 32'h7c000000),((LsuPlugin_pmaBuilder_io_addressBits & 32'hff000000) == 32'h7e000000)}}};
  assign _zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0_1 = _zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0[21];
  assign _zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0_2 = (_zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0[20] != early0_BranchPlugin_logic_alu_expectedMsb);
  assign _zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0_3 = (_zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0[19] != early0_BranchPlugin_logic_alu_expectedMsb);
  assign _zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0_4 = {(_zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0[18] != early0_BranchPlugin_logic_alu_expectedMsb),{(_zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0[17] != early0_BranchPlugin_logic_alu_expectedMsb),{(_zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0[16] != early0_BranchPlugin_logic_alu_expectedMsb),{(_zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0[15] != early0_BranchPlugin_logic_alu_expectedMsb),{(_zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0[14] != early0_BranchPlugin_logic_alu_expectedMsb),{(_zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0_5 != early0_BranchPlugin_logic_alu_expectedMsb),{_zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0_6,{_zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0_7,_zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0_8}}}}}}}};
  assign _zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0_5 = _zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0[13];
  assign _zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0_6 = (_zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0[12] != early0_BranchPlugin_logic_alu_expectedMsb);
  assign _zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0_7 = (_zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0[11] != early0_BranchPlugin_logic_alu_expectedMsb);
  assign _zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0_8 = {(_zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0[10] != early0_BranchPlugin_logic_alu_expectedMsb),{(_zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0[9] != early0_BranchPlugin_logic_alu_expectedMsb),{(_zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0[8] != early0_BranchPlugin_logic_alu_expectedMsb),{(_zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0[7] != early0_BranchPlugin_logic_alu_expectedMsb),{(_zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0[6] != early0_BranchPlugin_logic_alu_expectedMsb),{(_zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0_9 != early0_BranchPlugin_logic_alu_expectedMsb),{_zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0_10,{_zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0_11,_zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0_12}}}}}}}};
  assign _zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0_9 = _zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0[5];
  assign _zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0_10 = (_zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0[4] != early0_BranchPlugin_logic_alu_expectedMsb);
  assign _zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0_11 = (_zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0[3] != early0_BranchPlugin_logic_alu_expectedMsb);
  assign _zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0_12 = {(_zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0[2] != early0_BranchPlugin_logic_alu_expectedMsb),{(_zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0[1] != early0_BranchPlugin_logic_alu_expectedMsb),(_zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0[0] != early0_BranchPlugin_logic_alu_expectedMsb)}};
  assign _zz_decode_ctrls_1_down_RS1_ENABLE_0_1 = 32'h00005004;
  assign _zz_decode_ctrls_1_down_RS1_ENABLE_0_2 = 32'h00002050;
  assign _zz_decode_ctrls_1_down_RD_ENABLE_0_1 = 32'h00000050;
  assign _zz_decode_ctrls_1_down_RD_ENABLE_0_2 = (decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000000c);
  assign _zz_decode_ctrls_1_down_RD_ENABLE_0_3 = 32'h00000004;
  assign _zz_decode_ctrls_1_down_RD_ENABLE_0_4 = (decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000028);
  assign _zz_decode_ctrls_1_down_RD_ENABLE_0_5 = 32'h0;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0 = 32'h0000106f;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_1 = (decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000405f);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_2 = 32'h00000003;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_3 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000207f) == 32'h00002073);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_4 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000306f) == 32'h00001063);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_5 = {((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000407f) == 32'h00004063),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000207f) == 32'h00002013),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & _zz_decode_ctrls_1_down_Decode_LEGAL_0_6) == 32'h00000003),{(_zz_decode_ctrls_1_down_Decode_LEGAL_0_7 == _zz_decode_ctrls_1_down_Decode_LEGAL_0_8),{_zz_decode_ctrls_1_down_Decode_LEGAL_0_9,{_zz_decode_ctrls_1_down_Decode_LEGAL_0_10,_zz_decode_ctrls_1_down_Decode_LEGAL_0_11}}}}}};
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_6 = 32'h0000207f;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_7 = (decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000707b);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_8 = 32'h00000063;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_9 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000607f) == 32'h0000000f);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_10 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00007077) == 32'h00000013);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_11 = {((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h1800607f) == 32'h0000202f),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'he800607f) == 32'h0800202f),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & _zz_decode_ctrls_1_down_Decode_LEGAL_0_12) == 32'h00000033),{(_zz_decode_ctrls_1_down_Decode_LEGAL_0_13 == _zz_decode_ctrls_1_down_Decode_LEGAL_0_14),{_zz_decode_ctrls_1_down_Decode_LEGAL_0_15,{_zz_decode_ctrls_1_down_Decode_LEGAL_0_16,_zz_decode_ctrls_1_down_Decode_LEGAL_0_17}}}}}};
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_12 = 32'hfc00007f;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_13 = (decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hfe004077);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_14 = 32'h02004033;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_15 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hbc007077) == 32'h00005013);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_16 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hfc003077) == 32'h00001013);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_17 = {((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hbe007077) == 32'h00005033),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hfe003077) == 32'h02000033),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & _zz_decode_ctrls_1_down_Decode_LEGAL_0_18) == 32'h00001033),{(_zz_decode_ctrls_1_down_Decode_LEGAL_0_19 == _zz_decode_ctrls_1_down_Decode_LEGAL_0_20),{_zz_decode_ctrls_1_down_Decode_LEGAL_0_21,{_zz_decode_ctrls_1_down_Decode_LEGAL_0_22,_zz_decode_ctrls_1_down_Decode_LEGAL_0_23}}}}}};
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_18 = 32'hfe003077;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_19 = (decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hbe007077);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_20 = 32'h00000033;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_21 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hf9f0607f) == 32'h1000202f);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_22 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hfe007fff) == 32'h12000073);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_23 = {((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hffd07fff) == 32'h0000200f),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hffe07fff) == 32'h0000200f),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & _zz_decode_ctrls_1_down_Decode_LEGAL_0_24) == 32'h10200073),{(_zz_decode_ctrls_1_down_Decode_LEGAL_0_25 == _zz_decode_ctrls_1_down_Decode_LEGAL_0_26),(_zz_decode_ctrls_1_down_Decode_LEGAL_0_27 == _zz_decode_ctrls_1_down_Decode_LEGAL_0_28)}}}};
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_24 = 32'hdfffffff;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_25 = (decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hffefffff);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_26 = 32'h00000073;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_27 = (decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hffffffff);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_28 = 32'h10500073;
  assign _zz_CsrRamPlugin_csrMapper_ramAddress_1 = (_zz_CsrRamPlugin_csrMapper_ramAddress & 12'ha02);
  assign _zz_CsrRamPlugin_csrMapper_ramAddress_2 = 12'h202;
  assign _zz_CsrRamPlugin_csrMapper_ramAddress_3 = (_zz_CsrRamPlugin_csrMapper_ramAddress & 12'ha40);
  assign _zz_CsrRamPlugin_csrMapper_ramAddress_4 = 12'h200;
  assign _zz_CsrRamPlugin_csrMapper_ramAddress_5 = ((_zz_CsrRamPlugin_csrMapper_ramAddress & 12'ha02) == 12'h002);
  assign _zz_CsrRamPlugin_csrMapper_ramAddress_6 = ((_zz_CsrRamPlugin_csrMapper_ramAddress & _zz_CsrRamPlugin_csrMapper_ramAddress_7) == 12'h0);
  assign _zz_CsrRamPlugin_csrMapper_ramAddress_8 = ((_zz_CsrRamPlugin_csrMapper_ramAddress & _zz_CsrRamPlugin_csrMapper_ramAddress_9) == 12'h200);
  assign _zz_CsrRamPlugin_csrMapper_ramAddress_10 = ((_zz_CsrRamPlugin_csrMapper_ramAddress & 12'h806) == 12'h0);
  assign _zz_CsrRamPlugin_csrMapper_ramAddress_11 = ((_zz_CsrRamPlugin_csrMapper_ramAddress & _zz_CsrRamPlugin_csrMapper_ramAddress_12) == 12'h001);
  assign _zz_CsrRamPlugin_csrMapper_ramAddress_13 = ((_zz_CsrRamPlugin_csrMapper_ramAddress & _zz_CsrRamPlugin_csrMapper_ramAddress_14) == 12'h0);
  assign _zz_CsrRamPlugin_csrMapper_ramAddress_7 = 12'ha40;
  assign _zz_CsrRamPlugin_csrMapper_ramAddress_9 = 12'ha06;
  assign _zz_CsrRamPlugin_csrMapper_ramAddress_12 = 12'h003;
  assign _zz_CsrRamPlugin_csrMapper_ramAddress_14 = 12'h042;
  assign _zz_GSharePlugin_logic_onLearn_hash_1 = _zz_GSharePlugin_logic_onLearn_hash[6];
  assign _zz_GSharePlugin_logic_onLearn_hash_2 = _zz_GSharePlugin_logic_onLearn_hash[7];
  assign _zz_GSharePlugin_logic_onLearn_hash_3 = {_zz_GSharePlugin_logic_onLearn_hash[8],{_zz_GSharePlugin_logic_onLearn_hash[9],{_zz_GSharePlugin_logic_onLearn_hash[10],{_zz_GSharePlugin_logic_onLearn_hash[11],_zz_GSharePlugin_logic_onLearn_hash[12]}}}};
  assign _zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception = {TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_tval,TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_exception};
  assign _zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception_1 = {TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_tval,TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_exception};
  assign _zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception_2 = {TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_tval,TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_exception};
  assign _zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception_3 = {TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_tval,TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_exception};
  assign _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated = execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_physicalAddress;
  assign _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_1 = execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[11 : 0];
  assign _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_2 = execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_physicalAddress;
  assign _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_3 = execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[11 : 0];
  assign _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_4 = execute_ctrl3_down_MMU_L0_ENTRIES_lane0_2_physicalAddress;
  assign _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_5 = execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[11 : 0];
  assign _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_6 = execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_physicalAddress;
  assign _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_7 = execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[20 : 0];
  assign _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineTranslated = fetch_logic_ctrls_1_down_Fetch_WORD_PC[11 : 0];
  assign _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineTranslated_1 = fetch_logic_ctrls_1_down_Fetch_WORD_PC[11 : 0];
  assign _zz_fetch_logic_flushes_0_doIt = 1'b1;
  assign _zz_fetch_logic_flushes_0_doIt_1 = 1'b0;
  assign _zz_fetch_logic_flushes_0_doIt_2 = (1'b1 && BtbPlugin_logic_flushPort_payload_self);
  assign _zz_COMB_CSR_PmpPlugin_logic_allFilter = 12'h3bd;
  assign _zz_COMB_CSR_PmpPlugin_logic_allFilter_1 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h3bc);
  assign _zz_COMB_CSR_PmpPlugin_logic_allFilter_2 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h3bb);
  assign _zz_COMB_CSR_PmpPlugin_logic_allFilter_3 = {(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h3ba),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h3b9),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h3b8),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h3b7),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h3b6),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == _zz_COMB_CSR_PmpPlugin_logic_allFilter_4),{_zz_COMB_CSR_PmpPlugin_logic_allFilter_5,{_zz_COMB_CSR_PmpPlugin_logic_allFilter_6,_zz_COMB_CSR_PmpPlugin_logic_allFilter_7}}}}}}}};
  assign _zz_COMB_CSR_PmpPlugin_logic_allFilter_4 = 12'h3b5;
  assign _zz_COMB_CSR_PmpPlugin_logic_allFilter_5 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h3b4);
  assign _zz_COMB_CSR_PmpPlugin_logic_allFilter_6 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h3b3);
  assign _zz_COMB_CSR_PmpPlugin_logic_allFilter_7 = {(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h3b2),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h3b1),(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h3b0)}};
  assign _zz_COMB_CSR_UNAMED_1 = 12'h33d;
  assign _zz_COMB_CSR_UNAMED_1_1 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc1d);
  assign _zz_COMB_CSR_UNAMED_1_2 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb1d);
  assign _zz_COMB_CSR_UNAMED_1_3 = {(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h33c),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc1c),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb1c),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h33b),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc1b),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == _zz_COMB_CSR_UNAMED_1_4),{_zz_COMB_CSR_UNAMED_1_5,{_zz_COMB_CSR_UNAMED_1_6,_zz_COMB_CSR_UNAMED_1_7}}}}}}}};
  assign _zz_COMB_CSR_UNAMED_1_4 = 12'hb1b;
  assign _zz_COMB_CSR_UNAMED_1_5 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h33a);
  assign _zz_COMB_CSR_UNAMED_1_6 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc1a);
  assign _zz_COMB_CSR_UNAMED_1_7 = {(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb1a),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h339),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc19),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb19),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h338),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == _zz_COMB_CSR_UNAMED_1_8),{_zz_COMB_CSR_UNAMED_1_9,{_zz_COMB_CSR_UNAMED_1_10,_zz_COMB_CSR_UNAMED_1_11}}}}}}}};
  assign _zz_COMB_CSR_UNAMED_1_8 = 12'hc18;
  assign _zz_COMB_CSR_UNAMED_1_9 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb18);
  assign _zz_COMB_CSR_UNAMED_1_10 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h337);
  assign _zz_COMB_CSR_UNAMED_1_11 = {(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc17),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb17),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h336),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc16),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb16),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == _zz_COMB_CSR_UNAMED_1_12),{_zz_COMB_CSR_UNAMED_1_13,{_zz_COMB_CSR_UNAMED_1_14,_zz_COMB_CSR_UNAMED_1_15}}}}}}}};
  assign _zz_COMB_CSR_UNAMED_1_12 = 12'h335;
  assign _zz_COMB_CSR_UNAMED_1_13 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc15);
  assign _zz_COMB_CSR_UNAMED_1_14 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb15);
  assign _zz_COMB_CSR_UNAMED_1_15 = {(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h334),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc14),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb14),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h333),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc13),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == _zz_COMB_CSR_UNAMED_1_16),{_zz_COMB_CSR_UNAMED_1_17,{_zz_COMB_CSR_UNAMED_1_18,_zz_COMB_CSR_UNAMED_1_19}}}}}}}};
  assign _zz_COMB_CSR_UNAMED_1_16 = 12'hb13;
  assign _zz_COMB_CSR_UNAMED_1_17 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h332);
  assign _zz_COMB_CSR_UNAMED_1_18 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc12);
  assign _zz_COMB_CSR_UNAMED_1_19 = {(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb12),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h331),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc11),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb11),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h330),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == _zz_COMB_CSR_UNAMED_1_20),{_zz_COMB_CSR_UNAMED_1_21,{_zz_COMB_CSR_UNAMED_1_22,_zz_COMB_CSR_UNAMED_1_23}}}}}}}};
  assign _zz_COMB_CSR_UNAMED_1_20 = 12'hc10;
  assign _zz_COMB_CSR_UNAMED_1_21 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb10);
  assign _zz_COMB_CSR_UNAMED_1_22 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h32f);
  assign _zz_COMB_CSR_UNAMED_1_23 = {(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc0f),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb0f),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h32e),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc0e),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb0e),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == _zz_COMB_CSR_UNAMED_1_24),{_zz_COMB_CSR_UNAMED_1_25,{_zz_COMB_CSR_UNAMED_1_26,_zz_COMB_CSR_UNAMED_1_27}}}}}}}};
  assign _zz_COMB_CSR_UNAMED_1_24 = 12'h32d;
  assign _zz_COMB_CSR_UNAMED_1_25 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc0d);
  assign _zz_COMB_CSR_UNAMED_1_26 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb0d);
  assign _zz_COMB_CSR_UNAMED_1_27 = {(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h32c),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc0c),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb0c),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h32b),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc0b),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == _zz_COMB_CSR_UNAMED_1_28),{_zz_COMB_CSR_UNAMED_1_29,{_zz_COMB_CSR_UNAMED_1_30,_zz_COMB_CSR_UNAMED_1_31}}}}}}}};
  assign _zz_COMB_CSR_UNAMED_1_28 = 12'hb0b;
  assign _zz_COMB_CSR_UNAMED_1_29 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h32a);
  assign _zz_COMB_CSR_UNAMED_1_30 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc0a);
  assign _zz_COMB_CSR_UNAMED_1_31 = {(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb0a),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h329),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc09),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb09),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h328),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == _zz_COMB_CSR_UNAMED_1_32),{_zz_COMB_CSR_UNAMED_1_33,{_zz_COMB_CSR_UNAMED_1_34,_zz_COMB_CSR_UNAMED_1_35}}}}}}}};
  assign _zz_COMB_CSR_UNAMED_1_32 = 12'hc08;
  assign _zz_COMB_CSR_UNAMED_1_33 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb08);
  assign _zz_COMB_CSR_UNAMED_1_34 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h327);
  assign _zz_COMB_CSR_UNAMED_1_35 = {(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc07),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb07),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h326),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc06),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb06),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == _zz_COMB_CSR_UNAMED_1_36),{_zz_COMB_CSR_UNAMED_1_37,{_zz_COMB_CSR_UNAMED_1_38,_zz_COMB_CSR_UNAMED_1_39}}}}}}}};
  assign _zz_COMB_CSR_UNAMED_1_36 = 12'h325;
  assign _zz_COMB_CSR_UNAMED_1_37 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc05);
  assign _zz_COMB_CSR_UNAMED_1_38 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb05);
  assign _zz_COMB_CSR_UNAMED_1_39 = {(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h324),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc04),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb04),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h323),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc03),(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb03)}}}}};
  assign _zz_COMB_CSR_CsrRamPlugin_csrMapper_selFilter = 12'h143;
  assign _zz_COMB_CSR_CsrRamPlugin_csrMapper_selFilter_1 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h105);
  assign _zz_COMB_CSR_CsrRamPlugin_csrMapper_selFilter_2 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h340);
  assign _zz_COMB_CSR_CsrRamPlugin_csrMapper_selFilter_3 = {(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h341),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h343),(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h305)}};
  assign _zz_CsrAccessPlugin_logic_fsm_inject_implemented = COMB_CSR_3504;
  assign _zz_CsrAccessPlugin_logic_fsm_inject_implemented_1 = {COMB_CSR_324,{COMB_CSR_260,{COMB_CSR_778,{COMB_CSR_322,{COMB_CSR_774,{COMB_CSR_4016,{COMB_CSR_771,{COMB_CSR_770,{COMB_CSR_772,{COMB_CSR_836,{_zz_CsrAccessPlugin_logic_fsm_inject_implemented_2,_zz_CsrAccessPlugin_logic_fsm_inject_implemented_3}}}}}}}}}}};
  assign _zz_CsrAccessPlugin_logic_fsm_inject_implemented_2 = COMB_CSR_834;
  assign _zz_CsrAccessPlugin_logic_fsm_inject_implemented_3 = {COMB_CSR_769,{COMB_CSR_3860,{COMB_CSR_3859,{COMB_CSR_3858,{COMB_CSR_3857,{COMB_CSR_1954,{COMB_CSR_1953,{COMB_CSR_1952,{COMB_CSR_794,{COMB_CSR_PmpPlugin_logic_allFilter,{_zz_CsrAccessPlugin_logic_fsm_inject_implemented_4,_zz_CsrAccessPlugin_logic_fsm_inject_implemented_5}}}}}}}}}}};
  assign _zz_CsrAccessPlugin_logic_fsm_inject_implemented_4 = COMB_CSR_947;
  assign _zz_CsrAccessPlugin_logic_fsm_inject_implemented_5 = {COMB_CSR_946,{COMB_CSR_945,{COMB_CSR_928,{COMB_CSR_944,{COMB_CSR_384,{COMB_CSR_256,COMB_CSR_768}}}}}};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_32 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_33 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_38);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_43 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_44 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_48);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_53 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_54 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_59);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_64 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_65 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_70);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_75 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_76 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_81);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_86 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_87 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_92);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_97 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_98 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_103);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_108 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_109 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_114);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_119 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_120 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_125);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_128 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_129 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_132);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_133 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_134 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_139);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_143 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_144 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_149);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_154 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_155 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_160);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_164 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_165 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_170);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_175 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_176 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_181);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_186 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_187 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_192);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_197 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_198 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_203);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_208 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_209 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_214);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_219 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_220 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_224);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_228 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_229 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_234);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_239 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_240 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_245);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_249 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_250 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_255);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_260 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_261 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_266);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_271 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_272 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_277);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_282 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_283 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_288);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_291 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_292 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_297);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_302 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_303 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_308);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_313 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_314 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_317);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_33 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_34 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_36);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_38 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_39 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_41);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_44 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_45 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_46);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_48 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_49 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_51);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_54 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_55 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_57);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_59 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_60 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_62);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_65 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_66 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_68);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_70 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_71 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_73);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_76 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_77 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_79);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_81 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_82 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_84);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_87 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_88 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_90);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_92 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_93 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_95);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_98 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_99 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_101);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_103 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_104 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_106);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_109 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_110 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_112);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_114 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_115 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_117);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_120 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_121 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_123);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_125 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_126 | 64'h0);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_129 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_130 | 64'h0);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_132 = (64'h0 | ((when_CsrService_l232 && REG_CSR_769) ? 64'h8000000000141105 : 64'h0));
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_134 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_135 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_137);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_139 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_140 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_142);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_144 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_145 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_147);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_149 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_150 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_152);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_155 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_156 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_158);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_160 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_161 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_163);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_165 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_166 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_168);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_170 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_171 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_173);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_176 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_177 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_179);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_181 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_182 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_184);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_187 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_188 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_190);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_192 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_193 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_195);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_198 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_199 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_201);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_203 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_204 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_206);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_209 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_210 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_212);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_214 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_215 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_217);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_220 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_221 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_222);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_224 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_225 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_226);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_229 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_230 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_232);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_234 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_235 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_237);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_240 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_241 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_243);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_245 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_246 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_247);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_250 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_251 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_253);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_255 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_256 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_258);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_261 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_262 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_264);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_266 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_267 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_269);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_272 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_273 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_275);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_277 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_278 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_280);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_283 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_284 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_286);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_288 = (((when_CsrService_l232 && REG_CSR_3073) ? PrivilegedPlugin_logic_rdtime : 64'h0) | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_289);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_292 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_293 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_295);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_297 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_298 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_300);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_303 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_304 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_306);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_308 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_309 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_311);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_314 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_315 | (CsrRamPlugin_csrMapper_withRead ? CsrRamPlugin_csrMapper_read_data : 64'h0));
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_317 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_318 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_320);
  assign _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0 = 32'h00000010;
  assign _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0_1 = (execute_lane0_logic_decoding_decodingBits & 32'h00002020);
  assign _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0_2 = 32'h00002000;
  assign _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0_3 = ((execute_lane0_logic_decoding_decodingBits & 32'h08002000) == 32'h00002000);
  assign _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0_4 = 32'h00000018;
  assign _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0_5 = (execute_lane0_logic_decoding_decodingBits & 32'h00001008);
  assign _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0_6 = 32'h00001000;
  assign _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0_7 = ((execute_lane0_logic_decoding_decodingBits & 32'h10001010) == 32'h00001000);
  assign _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0_8 = ((execute_lane0_logic_decoding_decodingBits & 32'h08001010) == 32'h00001000);
  assign _zz__zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2 = 32'h02001000;
  assign _zz__zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_1 = 32'h10201000;
  assign _zz__zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_2 = (execute_lane0_logic_decoding_decodingBits & 32'h12400000);
  assign _zz__zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_3 = 32'h10000000;
  assign _zz__zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_4 = ((execute_lane0_logic_decoding_decodingBits & 32'h10100000) == 32'h00100000);
  assign _zz__zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_5 = ((execute_lane0_logic_decoding_decodingBits & 32'h12200000) == 32'h10000000);
  assign _zz_when_ExecuteLanePlugin_l306_2 = 1'b1;
  assign _zz_when_ExecuteLanePlugin_l306_2_1 = 1'b1;
  assign _zz_when_ExecuteLanePlugin_l306_2_2 = 1'b0;
  assign _zz_when_ExecuteLanePlugin_l306_2_3 = (1'b1 && early0_BranchPlugin_logic_flushPort_payload_self);
  assign BtbPlugin_logic_ras_mem_stack_spinal_port0 = BtbPlugin_logic_ras_mem_stack[BtbPlugin_logic_ras_ptr_pop_aheadValue];
  always @(posedge clk) begin
    if(_zz_3) begin
      BtbPlugin_logic_ras_mem_stack[BtbPlugin_logic_ras_write_payload_address] <= _zz_BtbPlugin_logic_ras_mem_stack_port;
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_banks_0_mem_spinal_port1 = {_zz_LsuL1Plugin_logic_banks_0_memsymbol_read_7, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_6, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_5, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_4, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_3, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_2, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_1, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read};
  end
  always @(posedge clk) begin
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[0] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol0[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[7 : 0];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[1] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol1[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[15 : 8];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[2] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol2[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[23 : 16];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[3] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol3[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[31 : 24];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[4] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol4[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[39 : 32];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[5] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol5[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[47 : 40];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[6] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol6[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[55 : 48];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[7] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol7[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[63 : 56];
    end
  end

  always @(posedge clk) begin
    if(LsuL1Plugin_logic_banks_0_read_cmd_valid) begin
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read <= LsuL1Plugin_logic_banks_0_mem_symbol0[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_1 <= LsuL1Plugin_logic_banks_0_mem_symbol1[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_2 <= LsuL1Plugin_logic_banks_0_mem_symbol2[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_3 <= LsuL1Plugin_logic_banks_0_mem_symbol3[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_4 <= LsuL1Plugin_logic_banks_0_mem_symbol4[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_5 <= LsuL1Plugin_logic_banks_0_mem_symbol5[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_6 <= LsuL1Plugin_logic_banks_0_mem_symbol6[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_7 <= LsuL1Plugin_logic_banks_0_mem_symbol7[LsuL1Plugin_logic_banks_0_read_cmd_payload];
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_banks_1_mem_spinal_port1 = {_zz_LsuL1Plugin_logic_banks_1_memsymbol_read_7, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_6, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_5, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_4, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_3, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_2, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_1, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read};
  end
  always @(posedge clk) begin
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[0] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol0[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[7 : 0];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[1] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol1[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[15 : 8];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[2] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol2[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[23 : 16];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[3] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol3[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[31 : 24];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[4] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol4[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[39 : 32];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[5] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol5[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[47 : 40];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[6] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol6[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[55 : 48];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[7] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol7[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[63 : 56];
    end
  end

  always @(posedge clk) begin
    if(LsuL1Plugin_logic_banks_1_read_cmd_valid) begin
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read <= LsuL1Plugin_logic_banks_1_mem_symbol0[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_1 <= LsuL1Plugin_logic_banks_1_mem_symbol1[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_2 <= LsuL1Plugin_logic_banks_1_mem_symbol2[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_3 <= LsuL1Plugin_logic_banks_1_mem_symbol3[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_4 <= LsuL1Plugin_logic_banks_1_mem_symbol4[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_5 <= LsuL1Plugin_logic_banks_1_mem_symbol5[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_6 <= LsuL1Plugin_logic_banks_1_mem_symbol6[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_7 <= LsuL1Plugin_logic_banks_1_mem_symbol7[LsuL1Plugin_logic_banks_1_read_cmd_payload];
    end
  end

  always @(posedge clk) begin
    if(_zz_LsuL1Plugin_logic_ways_0_mem_port_1) begin
      LsuL1Plugin_logic_ways_0_mem[LsuL1Plugin_logic_waysWrite_address] <= _zz_LsuL1Plugin_logic_ways_0_mem_port;
    end
  end

  always @(posedge clk) begin
    if(LsuL1Plugin_logic_ways_0_lsuRead_cmd_valid) begin
      LsuL1Plugin_logic_ways_0_mem_spinal_port1 <= LsuL1Plugin_logic_ways_0_mem[LsuL1Plugin_logic_ways_0_lsuRead_cmd_payload];
    end
  end

  always @(posedge clk) begin
    if(_zz_LsuL1Plugin_logic_ways_1_mem_port_1) begin
      LsuL1Plugin_logic_ways_1_mem[LsuL1Plugin_logic_waysWrite_address] <= _zz_LsuL1Plugin_logic_ways_1_mem_port;
    end
  end

  always @(posedge clk) begin
    if(LsuL1Plugin_logic_ways_1_lsuRead_cmd_valid) begin
      LsuL1Plugin_logic_ways_1_mem_spinal_port1 <= LsuL1Plugin_logic_ways_1_mem[LsuL1Plugin_logic_ways_1_lsuRead_cmd_payload];
    end
  end

  always @(posedge clk) begin
    if(_zz_9) begin
      LsuL1Plugin_logic_shared_mem[LsuL1Plugin_logic_shared_write_payload_address] <= _zz_LsuL1Plugin_logic_shared_mem_port;
    end
  end

  always @(posedge clk) begin
    if(LsuL1Plugin_logic_shared_lsuRead_cmd_valid) begin
      LsuL1Plugin_logic_shared_mem_spinal_port1 <= LsuL1Plugin_logic_shared_mem[LsuL1Plugin_logic_shared_lsuRead_cmd_payload];
    end
  end

  always @(posedge clk) begin
    if(_zz_8) begin
      LsuL1Plugin_logic_writeback_victimBuffer[_zz_LsuL1Plugin_logic_writeback_victimBuffer_port] <= LsuL1Plugin_logic_writeback_read_readedData;
    end
  end

  always @(posedge clk) begin
    if(LsuL1Plugin_logic_writeback_write_bufferRead_ready) begin
      LsuL1Plugin_logic_writeback_victimBuffer_spinal_port1 <= LsuL1Plugin_logic_writeback_victimBuffer[_zz_LsuL1Plugin_logic_writeback_write_word];
    end
  end

  always @(posedge clk) begin
    if(_zz_7) begin
      FetchL1Plugin_logic_banks_0_mem[FetchL1Plugin_logic_banks_0_write_payload_address] <= FetchL1Plugin_logic_banks_0_write_payload_data;
    end
  end

  always @(posedge clk) begin
    if(FetchL1Plugin_logic_banks_0_read_cmd_valid) begin
      FetchL1Plugin_logic_banks_0_mem_spinal_port1 <= FetchL1Plugin_logic_banks_0_mem[FetchL1Plugin_logic_banks_0_read_cmd_payload];
    end
  end

  always @(posedge clk) begin
    if(_zz_6) begin
      FetchL1Plugin_logic_banks_1_mem[FetchL1Plugin_logic_banks_1_write_payload_address] <= FetchL1Plugin_logic_banks_1_write_payload_data;
    end
  end

  always @(posedge clk) begin
    if(FetchL1Plugin_logic_banks_1_read_cmd_valid) begin
      FetchL1Plugin_logic_banks_1_mem_spinal_port1 <= FetchL1Plugin_logic_banks_1_mem[FetchL1Plugin_logic_banks_1_read_cmd_payload];
    end
  end

  always @(posedge clk) begin
    if(_zz_FetchL1Plugin_logic_ways_0_mem_port_1) begin
      FetchL1Plugin_logic_ways_0_mem[FetchL1Plugin_logic_waysWrite_address] <= _zz_FetchL1Plugin_logic_ways_0_mem_port;
    end
  end

  always @(posedge clk) begin
    if(FetchL1Plugin_logic_ways_0_read_cmd_valid) begin
      FetchL1Plugin_logic_ways_0_mem_spinal_port1 <= FetchL1Plugin_logic_ways_0_mem[FetchL1Plugin_logic_ways_0_read_cmd_payload];
    end
  end

  always @(posedge clk) begin
    if(_zz_FetchL1Plugin_logic_ways_1_mem_port_1) begin
      FetchL1Plugin_logic_ways_1_mem[FetchL1Plugin_logic_waysWrite_address] <= _zz_FetchL1Plugin_logic_ways_1_mem_port;
    end
  end

  always @(posedge clk) begin
    if(FetchL1Plugin_logic_ways_1_read_cmd_valid) begin
      FetchL1Plugin_logic_ways_1_mem_spinal_port1 <= FetchL1Plugin_logic_ways_1_mem[FetchL1Plugin_logic_ways_1_read_cmd_payload];
    end
  end

  always @(posedge clk) begin
    if(_zz_5) begin
      FetchL1Plugin_logic_plru_mem[FetchL1Plugin_logic_plru_write_payload_address] <= FetchL1Plugin_logic_plru_write_payload_data_0;
    end
  end

  always @(posedge clk) begin
    if(FetchL1Plugin_logic_plru_read_cmd_valid) begin
      FetchL1Plugin_logic_plru_mem_spinal_port1 <= FetchL1Plugin_logic_plru_mem[FetchL1Plugin_logic_plru_read_cmd_payload];
    end
  end

  always @(posedge clk) begin
    if(_zz_4) begin
      GSharePlugin_logic_mem_banks_0[GSharePlugin_logic_mem_writes_0_payload_address] <= _zz_GSharePlugin_logic_mem_banks_0_port;
    end
  end

  always @(posedge clk) begin
    if(fetch_logic_ctrls_0_down_isReady) begin
      GSharePlugin_logic_mem_banks_0_spinal_port1 <= GSharePlugin_logic_mem_banks_0[_zz_GSharePlugin_logic_readRsp_readed_0_0];
    end
  end

  always @(posedge clk) begin
    if(BtbPlugin_logic_memDp_wp_payload_mask[0] && BtbPlugin_logic_memDp_wp_valid) begin
      BtbPlugin_logic_mem[BtbPlugin_logic_memDp_wp_payload_address] <= _zz_BtbPlugin_logic_mem_port;
    end
  end

  always @(posedge clk) begin
    if(BtbPlugin_logic_memDp_rp_cmd_valid) begin
      BtbPlugin_logic_mem_spinal_port1 <= BtbPlugin_logic_mem[BtbPlugin_logic_memDp_rp_cmd_payload];
    end
  end

  always @(posedge clk) begin
    if(_zz_FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_0_port_1) begin
      FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_0[FetchL1Plugin_logic_translationStorage_logic_sl_0_write_address] <= _zz_FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_0_port;
    end
  end

  assign FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_0_spinal_port1 = FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_0[FetchL1Plugin_logic_translationPort_logic_read_0_readAddress];
  always @(posedge clk) begin
    if(_zz_FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_1_port_1) begin
      FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_1[FetchL1Plugin_logic_translationStorage_logic_sl_0_write_address] <= _zz_FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_1_port;
    end
  end

  assign FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_1_spinal_port1 = FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_1[FetchL1Plugin_logic_translationPort_logic_read_0_readAddress];
  always @(posedge clk) begin
    if(_zz_FetchL1Plugin_logic_translationStorage_logic_sl_1_ways_0_port_1) begin
      FetchL1Plugin_logic_translationStorage_logic_sl_1_ways_0[FetchL1Plugin_logic_translationStorage_logic_sl_1_write_address] <= _zz_FetchL1Plugin_logic_translationStorage_logic_sl_1_ways_0_port;
    end
  end

  assign FetchL1Plugin_logic_translationStorage_logic_sl_1_ways_0_spinal_port1 = FetchL1Plugin_logic_translationStorage_logic_sl_1_ways_0[FetchL1Plugin_logic_translationPort_logic_read_1_readAddress];
  always @(posedge clk) begin
    if(_zz_LsuPlugin_logic_translationStorage_logic_sl_0_ways_0_port_1) begin
      LsuPlugin_logic_translationStorage_logic_sl_0_ways_0[LsuPlugin_logic_translationStorage_logic_sl_0_write_address] <= _zz_LsuPlugin_logic_translationStorage_logic_sl_0_ways_0_port;
    end
  end

  assign LsuPlugin_logic_translationStorage_logic_sl_0_ways_0_spinal_port1 = LsuPlugin_logic_translationStorage_logic_sl_0_ways_0[LsuPlugin_logic_onAddress0_translationPort_logic_read_0_readAddress];
  always @(posedge clk) begin
    if(_zz_LsuPlugin_logic_translationStorage_logic_sl_0_ways_1_port_1) begin
      LsuPlugin_logic_translationStorage_logic_sl_0_ways_1[LsuPlugin_logic_translationStorage_logic_sl_0_write_address] <= _zz_LsuPlugin_logic_translationStorage_logic_sl_0_ways_1_port;
    end
  end

  assign LsuPlugin_logic_translationStorage_logic_sl_0_ways_1_spinal_port1 = LsuPlugin_logic_translationStorage_logic_sl_0_ways_1[LsuPlugin_logic_onAddress0_translationPort_logic_read_0_readAddress];
  always @(posedge clk) begin
    if(_zz_LsuPlugin_logic_translationStorage_logic_sl_0_ways_2_port_1) begin
      LsuPlugin_logic_translationStorage_logic_sl_0_ways_2[LsuPlugin_logic_translationStorage_logic_sl_0_write_address] <= _zz_LsuPlugin_logic_translationStorage_logic_sl_0_ways_2_port;
    end
  end

  assign LsuPlugin_logic_translationStorage_logic_sl_0_ways_2_spinal_port1 = LsuPlugin_logic_translationStorage_logic_sl_0_ways_2[LsuPlugin_logic_onAddress0_translationPort_logic_read_0_readAddress];
  always @(posedge clk) begin
    if(_zz_LsuPlugin_logic_translationStorage_logic_sl_1_ways_0_port_1) begin
      LsuPlugin_logic_translationStorage_logic_sl_1_ways_0[LsuPlugin_logic_translationStorage_logic_sl_1_write_address] <= _zz_LsuPlugin_logic_translationStorage_logic_sl_1_ways_0_port;
    end
  end

  assign LsuPlugin_logic_translationStorage_logic_sl_1_ways_0_spinal_port1 = LsuPlugin_logic_translationStorage_logic_sl_1_ways_0[LsuPlugin_logic_onAddress0_translationPort_logic_read_1_readAddress];
  always @(posedge clk) begin
    if(_zz_2) begin
      CsrRamPlugin_logic_mem[CsrRamPlugin_logic_writeLogic_port_payload_address] <= CsrRamPlugin_logic_writeLogic_port_payload_data;
    end
  end

  always @(posedge clk) begin
    if(CsrRamPlugin_logic_readLogic_port_cmd_valid) begin
      CsrRamPlugin_logic_mem_spinal_port1 <= CsrRamPlugin_logic_mem[CsrRamPlugin_logic_readLogic_port_cmd_payload];
    end
  end

  DivRadix early0_DivPlugin_logic_processing_div (
    .io_flush                  (execute_ctrl2_down_isReady                                       ), //i
    .io_cmd_valid              (early0_DivPlugin_logic_processing_div_io_cmd_valid               ), //i
    .io_cmd_ready              (early0_DivPlugin_logic_processing_div_io_cmd_ready               ), //o
    .io_cmd_payload_a          (early0_DivPlugin_logic_processing_a_delay_1[63:0]                ), //i
    .io_cmd_payload_b          (early0_DivPlugin_logic_processing_b_delay_1[63:0]                ), //i
    .io_cmd_payload_normalized (1'b0                                                             ), //i
    .io_cmd_payload_iterations (6'bxxxxxx                                                        ), //i
    .io_rsp_valid              (early0_DivPlugin_logic_processing_div_io_rsp_valid               ), //o
    .io_rsp_ready              (1'b0                                                             ), //i
    .io_rsp_payload_result     (early0_DivPlugin_logic_processing_div_io_rsp_payload_result[63:0]), //o
    .io_rsp_payload_remain     (early0_DivPlugin_logic_processing_div_io_rsp_payload_remain[63:0]), //o
    .clk                       (clk                                                              ), //i
    .reset                     (reset                                                            )  //i
  );
  StreamArbiter LsuPlugin_logic_flusher_arbiter (
    .io_inputs_0_valid (TrapPlugin_logic_lsuL1Invalidate_0_cmd_valid     ), //i
    .io_inputs_0_ready (LsuPlugin_logic_flusher_arbiter_io_inputs_0_ready), //o
    .io_output_valid   (LsuPlugin_logic_flusher_arbiter_io_output_valid  ), //o
    .io_output_ready   (LsuPlugin_logic_flusher_arbiter_io_output_ready  ), //i
    .io_chosenOH       (LsuPlugin_logic_flusher_arbiter_io_chosenOH      ), //o
    .clk               (clk                                              ), //i
    .reset             (reset                                            )  //i
  );
  StreamArbiter_1 LsuPlugin_logic_onAddress0_arbiter (
    .io_inputs_0_valid              (LsuPlugin_logic_onAddress0_ls_port_valid                          ), //i
    .io_inputs_0_ready              (LsuPlugin_logic_onAddress0_arbiter_io_inputs_0_ready              ), //o
    .io_inputs_0_payload_op         (LsuPlugin_logic_onAddress0_ls_port_payload_op[2:0]                ), //i
    .io_inputs_0_payload_address    (LsuPlugin_logic_onAddress0_ls_port_payload_address[38:0]          ), //i
    .io_inputs_0_payload_size       (LsuPlugin_logic_onAddress0_ls_port_payload_size[1:0]              ), //i
    .io_inputs_0_payload_load       (LsuPlugin_logic_onAddress0_ls_port_payload_load                   ), //i
    .io_inputs_0_payload_store      (LsuPlugin_logic_onAddress0_ls_port_payload_store                  ), //i
    .io_inputs_0_payload_atomic     (LsuPlugin_logic_onAddress0_ls_port_payload_atomic                 ), //i
    .io_inputs_0_payload_clean      (LsuPlugin_logic_onAddress0_ls_port_payload_clean                  ), //i
    .io_inputs_0_payload_invalidate (LsuPlugin_logic_onAddress0_ls_port_payload_invalidate             ), //i
    .io_inputs_0_payload_storeId    (LsuPlugin_logic_onAddress0_ls_port_payload_storeId[11:0]          ), //i
    .io_inputs_1_valid              (LsuPlugin_logic_onAddress0_access_port_valid                      ), //i
    .io_inputs_1_ready              (LsuPlugin_logic_onAddress0_arbiter_io_inputs_1_ready              ), //o
    .io_inputs_1_payload_op         (LsuPlugin_logic_onAddress0_access_port_payload_op[2:0]            ), //i
    .io_inputs_1_payload_address    (LsuPlugin_logic_onAddress0_access_port_payload_address[38:0]      ), //i
    .io_inputs_1_payload_size       (LsuPlugin_logic_onAddress0_access_port_payload_size[1:0]          ), //i
    .io_inputs_1_payload_load       (LsuPlugin_logic_onAddress0_access_port_payload_load               ), //i
    .io_inputs_1_payload_store      (LsuPlugin_logic_onAddress0_access_port_payload_store              ), //i
    .io_inputs_1_payload_atomic     (LsuPlugin_logic_onAddress0_access_port_payload_atomic             ), //i
    .io_inputs_1_payload_clean      (LsuPlugin_logic_onAddress0_access_port_payload_clean              ), //i
    .io_inputs_1_payload_invalidate (LsuPlugin_logic_onAddress0_access_port_payload_invalidate         ), //i
    .io_inputs_1_payload_storeId    (LsuPlugin_logic_onAddress0_access_port_payload_storeId[11:0]      ), //i
    .io_inputs_2_valid              (LsuPlugin_logic_onAddress0_flush_port_valid                       ), //i
    .io_inputs_2_ready              (LsuPlugin_logic_onAddress0_arbiter_io_inputs_2_ready              ), //o
    .io_inputs_2_payload_op         (LsuPlugin_logic_onAddress0_flush_port_payload_op[2:0]             ), //i
    .io_inputs_2_payload_address    (LsuPlugin_logic_onAddress0_flush_port_payload_address[38:0]       ), //i
    .io_inputs_2_payload_size       (LsuPlugin_logic_onAddress0_flush_port_payload_size[1:0]           ), //i
    .io_inputs_2_payload_load       (LsuPlugin_logic_onAddress0_flush_port_payload_load                ), //i
    .io_inputs_2_payload_store      (LsuPlugin_logic_onAddress0_flush_port_payload_store               ), //i
    .io_inputs_2_payload_atomic     (LsuPlugin_logic_onAddress0_flush_port_payload_atomic              ), //i
    .io_inputs_2_payload_clean      (LsuPlugin_logic_onAddress0_flush_port_payload_clean               ), //i
    .io_inputs_2_payload_invalidate (LsuPlugin_logic_onAddress0_flush_port_payload_invalidate          ), //i
    .io_inputs_2_payload_storeId    (LsuPlugin_logic_onAddress0_flush_port_payload_storeId[11:0]       ), //i
    .io_output_valid                (LsuPlugin_logic_onAddress0_arbiter_io_output_valid                ), //o
    .io_output_ready                (LsuPlugin_logic_onAddress0_arbiter_io_output_ready                ), //i
    .io_output_payload_op           (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_op[2:0]      ), //o
    .io_output_payload_address      (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_address[38:0]), //o
    .io_output_payload_size         (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_size[1:0]    ), //o
    .io_output_payload_load         (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_load         ), //o
    .io_output_payload_store        (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_store        ), //o
    .io_output_payload_atomic       (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_atomic       ), //o
    .io_output_payload_clean        (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_clean        ), //o
    .io_output_payload_invalidate   (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_invalidate   ), //o
    .io_output_payload_storeId      (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_storeId[11:0]), //o
    .io_chosen                      (LsuPlugin_logic_onAddress0_arbiter_io_chosen[1:0]                 ), //o
    .io_chosenOH                    (LsuPlugin_logic_onAddress0_arbiter_io_chosenOH[2:0]               ), //o
    .clk                            (clk                                                               ), //i
    .reset                          (reset                                                             )  //i
  );
  StreamArbiter_2 streamArbiter_5 (
    .io_inputs_0_valid                                     (LearnPlugin_logic_buffered_0_valid                                         ), //i
    .io_inputs_0_ready                                     (streamArbiter_5_io_inputs_0_ready                                          ), //o
    .io_inputs_0_payload_pcOnLastSlice                     (LearnPlugin_logic_buffered_0_payload_pcOnLastSlice[38:0]                   ), //i
    .io_inputs_0_payload_pcTarget                          (LearnPlugin_logic_buffered_0_payload_pcTarget[38:0]                        ), //i
    .io_inputs_0_payload_taken                             (LearnPlugin_logic_buffered_0_payload_taken                                 ), //i
    .io_inputs_0_payload_isBranch                          (LearnPlugin_logic_buffered_0_payload_isBranch                              ), //i
    .io_inputs_0_payload_isPush                            (LearnPlugin_logic_buffered_0_payload_isPush                                ), //i
    .io_inputs_0_payload_isPop                             (LearnPlugin_logic_buffered_0_payload_isPop                                 ), //i
    .io_inputs_0_payload_wasWrong                          (LearnPlugin_logic_buffered_0_payload_wasWrong                              ), //i
    .io_inputs_0_payload_badPredictedTarget                (LearnPlugin_logic_buffered_0_payload_badPredictedTarget                    ), //i
    .io_inputs_0_payload_history                           (LearnPlugin_logic_buffered_0_payload_history[11:0]                         ), //i
    .io_inputs_0_payload_uopId                             (LearnPlugin_logic_buffered_0_payload_uopId[15:0]                           ), //i
    .io_inputs_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 (LearnPlugin_logic_buffered_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_0[1:0]), //i
    .io_inputs_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_1 (LearnPlugin_logic_buffered_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_1[1:0]), //i
    .io_output_valid                                       (streamArbiter_5_io_output_valid                                            ), //o
    .io_output_ready                                       (LearnPlugin_logic_arbitrated_ready                                         ), //i
    .io_output_payload_pcOnLastSlice                       (streamArbiter_5_io_output_payload_pcOnLastSlice[38:0]                      ), //o
    .io_output_payload_pcTarget                            (streamArbiter_5_io_output_payload_pcTarget[38:0]                           ), //o
    .io_output_payload_taken                               (streamArbiter_5_io_output_payload_taken                                    ), //o
    .io_output_payload_isBranch                            (streamArbiter_5_io_output_payload_isBranch                                 ), //o
    .io_output_payload_isPush                              (streamArbiter_5_io_output_payload_isPush                                   ), //o
    .io_output_payload_isPop                               (streamArbiter_5_io_output_payload_isPop                                    ), //o
    .io_output_payload_wasWrong                            (streamArbiter_5_io_output_payload_wasWrong                                 ), //o
    .io_output_payload_badPredictedTarget                  (streamArbiter_5_io_output_payload_badPredictedTarget                       ), //o
    .io_output_payload_history                             (streamArbiter_5_io_output_payload_history[11:0]                            ), //o
    .io_output_payload_uopId                               (streamArbiter_5_io_output_payload_uopId[15:0]                              ), //o
    .io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_0   (streamArbiter_5_io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_0[1:0]   ), //o
    .io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_1   (streamArbiter_5_io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_1[1:0]   ), //o
    .io_chosenOH                                           (streamArbiter_5_io_chosenOH                                                ), //o
    .clk                                                   (clk                                                                        ), //i
    .reset                                                 (reset                                                                      )  //i
  );
  StreamArbiter_3 MmuPlugin_logic_refill_arbiter (
    .io_inputs_0_valid                 (TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_cmd_valid   ), //i
    .io_inputs_0_ready                 (MmuPlugin_logic_refill_arbiter_io_inputs_0_ready              ), //o
    .io_inputs_0_payload_address       (bits_address[38:0]                                            ), //i
    .io_inputs_0_payload_storageId     (bits_storageId                                                ), //i
    .io_inputs_0_payload_storageEnable (bits_storageEnable                                            ), //i
    .io_output_valid                   (MmuPlugin_logic_refill_arbiter_io_output_valid                ), //o
    .io_output_ready                   (MmuPlugin_logic_refill_arbiter_io_output_ready                ), //i
    .io_output_payload_address         (MmuPlugin_logic_refill_arbiter_io_output_payload_address[38:0]), //o
    .io_output_payload_storageId       (MmuPlugin_logic_refill_arbiter_io_output_payload_storageId    ), //o
    .io_output_payload_storageEnable   (MmuPlugin_logic_refill_arbiter_io_output_payload_storageEnable), //o
    .io_chosenOH                       (MmuPlugin_logic_refill_arbiter_io_chosenOH                    ), //o
    .clk                               (clk                                                           ), //i
    .reset                             (reset                                                         )  //i
  );
  StreamArbiter_4 MmuPlugin_logic_invalidate_arbiter (
    .io_inputs_0_valid (TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidate_cmd_valid), //i
    .io_inputs_0_ready (MmuPlugin_logic_invalidate_arbiter_io_inputs_0_ready           ), //o
    .io_output_valid   (MmuPlugin_logic_invalidate_arbiter_io_output_valid             ), //o
    .io_output_ready   (MmuPlugin_logic_invalidate_arbiter_io_output_ready             ), //i
    .io_chosenOH       (MmuPlugin_logic_invalidate_arbiter_io_chosenOH                 ), //o
    .clk               (clk                                                            ), //i
    .reset             (reset                                                          )  //i
  );
  RegFileMem integer_RegFilePlugin_logic_regfile_fpga (
    .io_writes_0_valid   (integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_valid       ), //i
    .io_writes_0_address (integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_address[4:0]), //i
    .io_writes_0_data    (integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_data[63:0]  ), //i
    .io_writes_0_uopId   (integer_RegFilePlugin_logic_writeMerges_0_bus_uopId[15:0]        ), //i
    .io_reads_0_valid    (execute_lane0_bypasser_integer_RS1_port_valid                    ), //i
    .io_reads_0_address  (execute_lane0_bypasser_integer_RS1_port_address[4:0]             ), //i
    .io_reads_0_data     (integer_RegFilePlugin_logic_regfile_fpga_io_reads_0_data[63:0]   ), //o
    .io_reads_1_valid    (execute_lane0_bypasser_integer_RS2_port_valid                    ), //i
    .io_reads_1_address  (execute_lane0_bypasser_integer_RS2_port_address[4:0]             ), //i
    .io_reads_1_data     (integer_RegFilePlugin_logic_regfile_fpga_io_reads_1_data[63:0]   ), //o
    .clk                 (clk                                                              ), //i
    .reset               (reset                                                            )  //i
  );
  always @(*) begin
    case(LsuL1Plugin_logic_writeback_read_slotReadLast_payload_way)
      1'b0 : _zz_LsuL1Plugin_logic_writeback_read_readedData = LsuL1Plugin_logic_banks_0_read_rsp;
      default : _zz_LsuL1Plugin_logic_writeback_read_readedData = LsuL1Plugin_logic_banks_1_read_rsp;
    endcase
  end

  always @(*) begin
    case(_zz_57)
      2'b00 : _zz_56 = 2'b00;
      2'b01 : _zz_56 = 2'b01;
      2'b10 : _zz_56 = 2'b01;
      default : _zz_56 = 2'b10;
    endcase
  end

  always @(*) begin
    case(_zz_59)
      3'b000 : _zz_58 = 2'b00;
      3'b001 : _zz_58 = 2'b01;
      3'b010 : _zz_58 = 2'b01;
      3'b011 : _zz_58 = 2'b10;
      3'b100 : _zz_58 = 2'b01;
      3'b101 : _zz_58 = 2'b10;
      3'b110 : _zz_58 = 2'b10;
      default : _zz_58 = 2'b11;
    endcase
  end

  always @(*) begin
    case(LsuL1Plugin_logic_lsu_ctrl_needFlushSel)
      1'b0 : begin
        _zz__zz_LsuL1Plugin_logic_waysWrite_tag_address = execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_address;
        _zz_LsuL1Plugin_logic_waysWrite_tag_fault_1 = execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault;
      end
      default : begin
        _zz__zz_LsuL1Plugin_logic_waysWrite_tag_address = execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_address;
        _zz_LsuL1Plugin_logic_waysWrite_tag_fault_1 = execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault;
      end
    endcase
  end

  always @(*) begin
    case(LsuL1Plugin_logic_lsu_ctrl_targetWay)
      1'b0 : _zz_LsuL1Plugin_logic_writeback_push_payload_address = execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_address;
      default : _zz_LsuL1Plugin_logic_writeback_push_payload_address = execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_address;
    endcase
  end

  always @(*) begin
    case(_zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_0_1)
      1'b0 : _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_0 = fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_WORDS_0[31 : 0];
      default : _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_0 = fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_WORDS_0[63 : 32];
    endcase
  end

  always @(*) begin
    case(_zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_1_1)
      1'b0 : _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_1 = fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_WORDS_1[31 : 0];
      default : _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_1 = fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_WORDS_1[63 : 32];
    endcase
  end

  always @(*) begin
    case(_zz_PerformanceCounterPlugin_logic_commitCount_1)
      1'b0 : _zz_PerformanceCounterPlugin_logic_commitCount = 1'b0;
      default : _zz_PerformanceCounterPlugin_logic_commitCount = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_LsuPlugin_logic_onCtrl_loadData_shifted_1)
      3'b000 : _zz_LsuPlugin_logic_onCtrl_loadData_shifted = LsuPlugin_logic_onCtrl_loadData_splitted_0;
      3'b001 : _zz_LsuPlugin_logic_onCtrl_loadData_shifted = LsuPlugin_logic_onCtrl_loadData_splitted_1;
      3'b010 : _zz_LsuPlugin_logic_onCtrl_loadData_shifted = LsuPlugin_logic_onCtrl_loadData_splitted_2;
      3'b011 : _zz_LsuPlugin_logic_onCtrl_loadData_shifted = LsuPlugin_logic_onCtrl_loadData_splitted_3;
      3'b100 : _zz_LsuPlugin_logic_onCtrl_loadData_shifted = LsuPlugin_logic_onCtrl_loadData_splitted_4;
      3'b101 : _zz_LsuPlugin_logic_onCtrl_loadData_shifted = LsuPlugin_logic_onCtrl_loadData_splitted_5;
      3'b110 : _zz_LsuPlugin_logic_onCtrl_loadData_shifted = LsuPlugin_logic_onCtrl_loadData_splitted_6;
      default : _zz_LsuPlugin_logic_onCtrl_loadData_shifted = LsuPlugin_logic_onCtrl_loadData_splitted_7;
    endcase
  end

  always @(*) begin
    case(_zz_LsuPlugin_logic_onCtrl_loadData_shifted_3)
      2'b00 : _zz_LsuPlugin_logic_onCtrl_loadData_shifted_2 = LsuPlugin_logic_onCtrl_loadData_splitted_1;
      2'b01 : _zz_LsuPlugin_logic_onCtrl_loadData_shifted_2 = LsuPlugin_logic_onCtrl_loadData_splitted_3;
      2'b10 : _zz_LsuPlugin_logic_onCtrl_loadData_shifted_2 = LsuPlugin_logic_onCtrl_loadData_splitted_5;
      default : _zz_LsuPlugin_logic_onCtrl_loadData_shifted_2 = LsuPlugin_logic_onCtrl_loadData_splitted_7;
    endcase
  end

  always @(*) begin
    case(_zz_LsuPlugin_logic_onCtrl_loadData_shifted_5)
      1'b0 : _zz_LsuPlugin_logic_onCtrl_loadData_shifted_4 = LsuPlugin_logic_onCtrl_loadData_splitted_2;
      default : _zz_LsuPlugin_logic_onCtrl_loadData_shifted_4 = LsuPlugin_logic_onCtrl_loadData_splitted_6;
    endcase
  end

  always @(*) begin
    case(_zz_LsuPlugin_logic_onCtrl_loadData_shifted_7)
      1'b0 : _zz_LsuPlugin_logic_onCtrl_loadData_shifted_6 = LsuPlugin_logic_onCtrl_loadData_splitted_3;
      default : _zz_LsuPlugin_logic_onCtrl_loadData_shifted_6 = LsuPlugin_logic_onCtrl_loadData_splitted_7;
    endcase
  end

  always @(*) begin
    case(_zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK_1)
      1'b0 : _zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK = AlignerPlugin_logic_maskGen_frontMasks_0;
      default : _zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK = AlignerPlugin_logic_maskGen_frontMasks_1;
    endcase
  end

  always @(*) begin
    case(fetch_logic_ctrls_2_down_Prediction_WORD_JUMP_SLICE)
      1'b0 : _zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK_2 = AlignerPlugin_logic_maskGen_backMasks_0;
      default : _zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK_2 = AlignerPlugin_logic_maskGen_backMasks_1;
    endcase
  end

  always @(*) begin
    case(_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_24)
      2'b00 : _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_23 = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_18;
      2'b01 : _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_23 = (_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_18 | 32'h40000000);
      2'b10 : _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_23 = {{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_5,_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst},3'b111},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst},7'h13};
      default : _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_23 = ({{{{{7'h0,_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_1},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_25},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst},(AlignerPlugin_logic_extractors_0_ctx_instruction[12] ? 7'h3b : 7'h33)} | ((AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 5] == 2'b00) ? 32'h40000000 : 32'h0));
    endcase
  end

  always @(*) begin
    case(_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_26)
      3'b000 : _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_25 = 3'b000;
      3'b001 : _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_25 = 3'b100;
      3'b010 : _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_25 = 3'b110;
      3'b011 : _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_25 = 3'b111;
      3'b100 : _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_25 = 3'b000;
      3'b101 : _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_25 = 3'b000;
      3'b110 : _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_25 = 3'b010;
      default : _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_25 = 3'b011;
    endcase
  end

  always @(*) begin
    case(_zz_PerformanceCounterPlugin_logic_events_sums_0_2)
      1'b0 : _zz_PerformanceCounterPlugin_logic_events_sums_0_1 = 1'b0;
      default : _zz_PerformanceCounterPlugin_logic_events_sums_0_1 = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_PerformanceCounterPlugin_logic_events_sums_1_2)
      1'b0 : _zz_PerformanceCounterPlugin_logic_events_sums_1_1 = 1'b0;
      default : _zz_PerformanceCounterPlugin_logic_events_sums_1_1 = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_PerformanceCounterPlugin_logic_events_sums_2_2)
      1'b0 : _zz_PerformanceCounterPlugin_logic_events_sums_2_1 = 1'b0;
      default : _zz_PerformanceCounterPlugin_logic_events_sums_2_1 = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_PerformanceCounterPlugin_logic_events_sums_3_2)
      1'b0 : _zz_PerformanceCounterPlugin_logic_events_sums_3_1 = 1'b0;
      default : _zz_PerformanceCounterPlugin_logic_events_sums_3_1 = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_PerformanceCounterPlugin_logic_events_sums_4_2)
      1'b0 : _zz_PerformanceCounterPlugin_logic_events_sums_4_1 = 1'b0;
      default : _zz_PerformanceCounterPlugin_logic_events_sums_4_1 = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_PerformanceCounterPlugin_logic_events_sums_5_2)
      1'b0 : _zz_PerformanceCounterPlugin_logic_events_sums_5_1 = 1'b0;
      default : _zz_PerformanceCounterPlugin_logic_events_sums_5_1 = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_PerformanceCounterPlugin_logic_events_sums_6_2)
      1'b0 : _zz_PerformanceCounterPlugin_logic_events_sums_6_1 = 1'b0;
      default : _zz_PerformanceCounterPlugin_logic_events_sums_6_1 = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_PerformanceCounterPlugin_logic_events_sums_7_2)
      1'b0 : _zz_PerformanceCounterPlugin_logic_events_sums_7_1 = 1'b0;
      default : _zz_PerformanceCounterPlugin_logic_events_sums_7_1 = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_PerformanceCounterPlugin_logic_events_sums_8_2)
      1'b0 : _zz_PerformanceCounterPlugin_logic_events_sums_8_1 = 1'b0;
      default : _zz_PerformanceCounterPlugin_logic_events_sums_8_1 = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_PerformanceCounterPlugin_logic_events_sums_9_2)
      1'b0 : _zz_PerformanceCounterPlugin_logic_events_sums_9_1 = 1'b0;
      default : _zz_PerformanceCounterPlugin_logic_events_sums_9_1 = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_PerformanceCounterPlugin_logic_events_sums_10_2)
      1'b0 : _zz_PerformanceCounterPlugin_logic_events_sums_10_1 = 1'b0;
      default : _zz_PerformanceCounterPlugin_logic_events_sums_10_1 = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_PerformanceCounterPlugin_logic_events_sums_11_2)
      1'b0 : _zz_PerformanceCounterPlugin_logic_events_sums_11_1 = 1'b0;
      default : _zz_PerformanceCounterPlugin_logic_events_sums_11_1 = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_PerformanceCounterPlugin_logic_events_sums_12_2)
      1'b0 : _zz_PerformanceCounterPlugin_logic_events_sums_12_1 = 1'b0;
      default : _zz_PerformanceCounterPlugin_logic_events_sums_12_1 = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_PerformanceCounterPlugin_logic_events_sums_13_2)
      1'b0 : _zz_PerformanceCounterPlugin_logic_events_sums_13_1 = 1'b0;
      default : _zz_PerformanceCounterPlugin_logic_events_sums_13_1 = 1'b1;
    endcase
  end

  always @(*) begin
    case(CsrRamPlugin_logic_readLogic_sel)
      2'b00 : _zz_CsrRamPlugin_logic_readLogic_port_cmd_payload = PerformanceCounterPlugin_logic_readPort_address;
      2'b01 : _zz_CsrRamPlugin_logic_readLogic_port_cmd_payload = TrapPlugin_logic_harts_0_crsPorts_read_address;
      default : _zz_CsrRamPlugin_logic_readLogic_port_cmd_payload = CsrRamPlugin_csrMapper_read_address;
    endcase
  end

  always @(*) begin
    case(_zz_WhiteboxerPlugin_logic_perf_candidatesCount_1)
      1'b0 : _zz_WhiteboxerPlugin_logic_perf_candidatesCount = 1'b0;
      default : _zz_WhiteboxerPlugin_logic_perf_candidatesCount = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_WhiteboxerPlugin_logic_perf_dispatchFeedCount_1)
      1'b0 : _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCount = 1'b0;
      default : _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCount = 1'b1;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(execute_ctrl2_up_early0_EnvPlugin_OP_lane0)
      EnvPluginOp_ECALL : execute_ctrl2_up_early0_EnvPlugin_OP_lane0_string = "ECALL     ";
      EnvPluginOp_EBREAK : execute_ctrl2_up_early0_EnvPlugin_OP_lane0_string = "EBREAK    ";
      EnvPluginOp_PRIV_RET : execute_ctrl2_up_early0_EnvPlugin_OP_lane0_string = "PRIV_RET  ";
      EnvPluginOp_FENCE_I : execute_ctrl2_up_early0_EnvPlugin_OP_lane0_string = "FENCE_I   ";
      EnvPluginOp_SFENCE_VMA : execute_ctrl2_up_early0_EnvPlugin_OP_lane0_string = "SFENCE_VMA";
      EnvPluginOp_WFI : execute_ctrl2_up_early0_EnvPlugin_OP_lane0_string = "WFI       ";
      default : execute_ctrl2_up_early0_EnvPlugin_OP_lane0_string = "??????????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane0)
      BranchPlugin_BranchCtrlEnum_B : execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane0_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane0_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane0_string = "JALR";
      default : execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane0_string = "????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl2_up_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : execute_ctrl2_up_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : execute_ctrl2_up_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : execute_ctrl2_up_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : execute_ctrl2_up_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "ZERO ";
      default : execute_ctrl2_up_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "?????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl1_down_early0_EnvPlugin_OP_lane0)
      EnvPluginOp_ECALL : execute_ctrl1_down_early0_EnvPlugin_OP_lane0_string = "ECALL     ";
      EnvPluginOp_EBREAK : execute_ctrl1_down_early0_EnvPlugin_OP_lane0_string = "EBREAK    ";
      EnvPluginOp_PRIV_RET : execute_ctrl1_down_early0_EnvPlugin_OP_lane0_string = "PRIV_RET  ";
      EnvPluginOp_FENCE_I : execute_ctrl1_down_early0_EnvPlugin_OP_lane0_string = "FENCE_I   ";
      EnvPluginOp_SFENCE_VMA : execute_ctrl1_down_early0_EnvPlugin_OP_lane0_string = "SFENCE_VMA";
      EnvPluginOp_WFI : execute_ctrl1_down_early0_EnvPlugin_OP_lane0_string = "WFI       ";
      default : execute_ctrl1_down_early0_EnvPlugin_OP_lane0_string = "??????????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0)
      BranchPlugin_BranchCtrlEnum_B : execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_string = "JALR";
      default : execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_string = "????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "ZERO ";
      default : execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "?????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0)
      BranchPlugin_BranchCtrlEnum_B : execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0_string = "JALR";
      default : execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0_string = "????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl2_down_early0_EnvPlugin_OP_lane0)
      EnvPluginOp_ECALL : execute_ctrl2_down_early0_EnvPlugin_OP_lane0_string = "ECALL     ";
      EnvPluginOp_EBREAK : execute_ctrl2_down_early0_EnvPlugin_OP_lane0_string = "EBREAK    ";
      EnvPluginOp_PRIV_RET : execute_ctrl2_down_early0_EnvPlugin_OP_lane0_string = "PRIV_RET  ";
      EnvPluginOp_FENCE_I : execute_ctrl2_down_early0_EnvPlugin_OP_lane0_string = "FENCE_I   ";
      EnvPluginOp_SFENCE_VMA : execute_ctrl2_down_early0_EnvPlugin_OP_lane0_string = "SFENCE_VMA";
      EnvPluginOp_WFI : execute_ctrl2_down_early0_EnvPlugin_OP_lane0_string = "WFI       ";
      default : execute_ctrl2_down_early0_EnvPlugin_OP_lane0_string = "??????????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl2_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : execute_ctrl2_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : execute_ctrl2_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : execute_ctrl2_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : execute_ctrl2_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "ZERO ";
      default : execute_ctrl2_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "?????";
    endcase
  end
  always @(*) begin
    case(LsuPlugin_logic_onAddress0_ls_port_payload_op)
      LsuL1CmdOpcode_LSU : LsuPlugin_logic_onAddress0_ls_port_payload_op_string = "LSU         ";
      LsuL1CmdOpcode_ACCESS_1 : LsuPlugin_logic_onAddress0_ls_port_payload_op_string = "ACCESS_1    ";
      LsuL1CmdOpcode_STORE_BUFFER : LsuPlugin_logic_onAddress0_ls_port_payload_op_string = "STORE_BUFFER";
      LsuL1CmdOpcode_FLUSH : LsuPlugin_logic_onAddress0_ls_port_payload_op_string = "FLUSH       ";
      LsuL1CmdOpcode_PREFETCH : LsuPlugin_logic_onAddress0_ls_port_payload_op_string = "PREFETCH    ";
      default : LsuPlugin_logic_onAddress0_ls_port_payload_op_string = "????????????";
    endcase
  end
  always @(*) begin
    case(LsuPlugin_logic_onAddress0_access_port_payload_op)
      LsuL1CmdOpcode_LSU : LsuPlugin_logic_onAddress0_access_port_payload_op_string = "LSU         ";
      LsuL1CmdOpcode_ACCESS_1 : LsuPlugin_logic_onAddress0_access_port_payload_op_string = "ACCESS_1    ";
      LsuL1CmdOpcode_STORE_BUFFER : LsuPlugin_logic_onAddress0_access_port_payload_op_string = "STORE_BUFFER";
      LsuL1CmdOpcode_FLUSH : LsuPlugin_logic_onAddress0_access_port_payload_op_string = "FLUSH       ";
      LsuL1CmdOpcode_PREFETCH : LsuPlugin_logic_onAddress0_access_port_payload_op_string = "PREFETCH    ";
      default : LsuPlugin_logic_onAddress0_access_port_payload_op_string = "????????????";
    endcase
  end
  always @(*) begin
    case(LsuPlugin_logic_onAddress0_flush_port_payload_op)
      LsuL1CmdOpcode_LSU : LsuPlugin_logic_onAddress0_flush_port_payload_op_string = "LSU         ";
      LsuL1CmdOpcode_ACCESS_1 : LsuPlugin_logic_onAddress0_flush_port_payload_op_string = "ACCESS_1    ";
      LsuL1CmdOpcode_STORE_BUFFER : LsuPlugin_logic_onAddress0_flush_port_payload_op_string = "STORE_BUFFER";
      LsuL1CmdOpcode_FLUSH : LsuPlugin_logic_onAddress0_flush_port_payload_op_string = "FLUSH       ";
      LsuL1CmdOpcode_PREFETCH : LsuPlugin_logic_onAddress0_flush_port_payload_op_string = "PREFETCH    ";
      default : LsuPlugin_logic_onAddress0_flush_port_payload_op_string = "????????????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "ZERO ";
      default : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1_string = "ZERO ";
      default : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2_string = "ZERO ";
      default : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0)
      BranchPlugin_BranchCtrlEnum_B : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_string = "JALR";
      default : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_1)
      BranchPlugin_BranchCtrlEnum_B : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_1_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_1_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_1_string = "JALR";
      default : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_1_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_2)
      BranchPlugin_BranchCtrlEnum_B : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_2_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_2_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_2_string = "JALR";
      default : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_2_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1)
      EnvPluginOp_ECALL : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1_string = "ECALL     ";
      EnvPluginOp_EBREAK : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1_string = "EBREAK    ";
      EnvPluginOp_PRIV_RET : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1_string = "PRIV_RET  ";
      EnvPluginOp_FENCE_I : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1_string = "FENCE_I   ";
      EnvPluginOp_SFENCE_VMA : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1_string = "SFENCE_VMA";
      EnvPluginOp_WFI : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1_string = "WFI       ";
      default : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1_string = "??????????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2)
      EnvPluginOp_ECALL : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_string = "ECALL     ";
      EnvPluginOp_EBREAK : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_string = "EBREAK    ";
      EnvPluginOp_PRIV_RET : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_string = "PRIV_RET  ";
      EnvPluginOp_FENCE_I : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_string = "FENCE_I   ";
      EnvPluginOp_SFENCE_VMA : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_string = "SFENCE_VMA";
      EnvPluginOp_WFI : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_string = "WFI       ";
      default : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_string = "??????????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_3)
      EnvPluginOp_ECALL : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_3_string = "ECALL     ";
      EnvPluginOp_EBREAK : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_3_string = "EBREAK    ";
      EnvPluginOp_PRIV_RET : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_3_string = "PRIV_RET  ";
      EnvPluginOp_FENCE_I : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_3_string = "FENCE_I   ";
      EnvPluginOp_SFENCE_VMA : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_3_string = "SFENCE_VMA";
      EnvPluginOp_WFI : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_3_string = "WFI       ";
      default : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_3_string = "??????????";
    endcase
  end
  always @(*) begin
    case(LsuPlugin_logic_flusher_stateReg)
      LsuPlugin_logic_flusher_IDLE : LsuPlugin_logic_flusher_stateReg_string = "IDLE      ";
      LsuPlugin_logic_flusher_CMD : LsuPlugin_logic_flusher_stateReg_string = "CMD       ";
      LsuPlugin_logic_flusher_COMPLETION : LsuPlugin_logic_flusher_stateReg_string = "COMPLETION";
      default : LsuPlugin_logic_flusher_stateReg_string = "??????????";
    endcase
  end
  always @(*) begin
    case(LsuPlugin_logic_flusher_stateNext)
      LsuPlugin_logic_flusher_IDLE : LsuPlugin_logic_flusher_stateNext_string = "IDLE      ";
      LsuPlugin_logic_flusher_CMD : LsuPlugin_logic_flusher_stateNext_string = "CMD       ";
      LsuPlugin_logic_flusher_COMPLETION : LsuPlugin_logic_flusher_stateNext_string = "COMPLETION";
      default : LsuPlugin_logic_flusher_stateNext_string = "??????????";
    endcase
  end
  always @(*) begin
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RESET : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "RESET      ";
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "RUNNING    ";
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "COMPUTE    ";
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "TRAP_EPC   ";
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "TRAP_TVAL  ";
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "TRAP_TVEC  ";
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_WAIT : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "TRAP_WAIT  ";
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "TRAP_APPLY ";
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "XRET_EPC   ";
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "XRET_APPLY ";
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "ATS_RSP    ";
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "JUMP       ";
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "LSU_FLUSH  ";
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "FETCH_FLUSH";
      default : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "???????????";
    endcase
  end
  always @(*) begin
    case(TrapPlugin_logic_harts_0_trap_fsm_stateNext)
      TrapPlugin_logic_harts_0_trap_fsm_RESET : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "RESET      ";
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "RUNNING    ";
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "COMPUTE    ";
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "TRAP_EPC   ";
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "TRAP_TVAL  ";
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "TRAP_TVEC  ";
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_WAIT : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "TRAP_WAIT  ";
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "TRAP_APPLY ";
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "XRET_EPC   ";
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "XRET_APPLY ";
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "ATS_RSP    ";
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "JUMP       ";
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "LSU_FLUSH  ";
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "FETCH_FLUSH";
      default : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "???????????";
    endcase
  end
  always @(*) begin
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_BOOT : MmuPlugin_logic_refill_stateReg_string = "BOOT  ";
      MmuPlugin_logic_refill_IDLE : MmuPlugin_logic_refill_stateReg_string = "IDLE  ";
      MmuPlugin_logic_refill_CMD_0 : MmuPlugin_logic_refill_stateReg_string = "CMD_0 ";
      MmuPlugin_logic_refill_CMD_1 : MmuPlugin_logic_refill_stateReg_string = "CMD_1 ";
      MmuPlugin_logic_refill_CMD_2 : MmuPlugin_logic_refill_stateReg_string = "CMD_2 ";
      MmuPlugin_logic_refill_RSP_0 : MmuPlugin_logic_refill_stateReg_string = "RSP_0 ";
      MmuPlugin_logic_refill_RSP_1 : MmuPlugin_logic_refill_stateReg_string = "RSP_1 ";
      MmuPlugin_logic_refill_RSP_2 : MmuPlugin_logic_refill_stateReg_string = "RSP_2 ";
      MmuPlugin_logic_refill_DONE_0 : MmuPlugin_logic_refill_stateReg_string = "DONE_0";
      MmuPlugin_logic_refill_DONE_1 : MmuPlugin_logic_refill_stateReg_string = "DONE_1";
      MmuPlugin_logic_refill_DONE_2 : MmuPlugin_logic_refill_stateReg_string = "DONE_2";
      default : MmuPlugin_logic_refill_stateReg_string = "??????";
    endcase
  end
  always @(*) begin
    case(MmuPlugin_logic_refill_stateNext)
      MmuPlugin_logic_refill_BOOT : MmuPlugin_logic_refill_stateNext_string = "BOOT  ";
      MmuPlugin_logic_refill_IDLE : MmuPlugin_logic_refill_stateNext_string = "IDLE  ";
      MmuPlugin_logic_refill_CMD_0 : MmuPlugin_logic_refill_stateNext_string = "CMD_0 ";
      MmuPlugin_logic_refill_CMD_1 : MmuPlugin_logic_refill_stateNext_string = "CMD_1 ";
      MmuPlugin_logic_refill_CMD_2 : MmuPlugin_logic_refill_stateNext_string = "CMD_2 ";
      MmuPlugin_logic_refill_RSP_0 : MmuPlugin_logic_refill_stateNext_string = "RSP_0 ";
      MmuPlugin_logic_refill_RSP_1 : MmuPlugin_logic_refill_stateNext_string = "RSP_1 ";
      MmuPlugin_logic_refill_RSP_2 : MmuPlugin_logic_refill_stateNext_string = "RSP_2 ";
      MmuPlugin_logic_refill_DONE_0 : MmuPlugin_logic_refill_stateNext_string = "DONE_0";
      MmuPlugin_logic_refill_DONE_1 : MmuPlugin_logic_refill_stateNext_string = "DONE_1";
      MmuPlugin_logic_refill_DONE_2 : MmuPlugin_logic_refill_stateNext_string = "DONE_2";
      default : MmuPlugin_logic_refill_stateNext_string = "??????";
    endcase
  end
  always @(*) begin
    case(PerformanceCounterPlugin_logic_fsm_stateReg)
      PerformanceCounterPlugin_logic_fsm_BOOT : PerformanceCounterPlugin_logic_fsm_stateReg_string = "BOOT     ";
      PerformanceCounterPlugin_logic_fsm_IDLE : PerformanceCounterPlugin_logic_fsm_stateReg_string = "IDLE     ";
      PerformanceCounterPlugin_logic_fsm_READ_LOW : PerformanceCounterPlugin_logic_fsm_stateReg_string = "READ_LOW ";
      PerformanceCounterPlugin_logic_fsm_CALC_LOW : PerformanceCounterPlugin_logic_fsm_stateReg_string = "CALC_LOW ";
      PerformanceCounterPlugin_logic_fsm_CSR_WRITE : PerformanceCounterPlugin_logic_fsm_stateReg_string = "CSR_WRITE";
      default : PerformanceCounterPlugin_logic_fsm_stateReg_string = "?????????";
    endcase
  end
  always @(*) begin
    case(PerformanceCounterPlugin_logic_fsm_stateNext)
      PerformanceCounterPlugin_logic_fsm_BOOT : PerformanceCounterPlugin_logic_fsm_stateNext_string = "BOOT     ";
      PerformanceCounterPlugin_logic_fsm_IDLE : PerformanceCounterPlugin_logic_fsm_stateNext_string = "IDLE     ";
      PerformanceCounterPlugin_logic_fsm_READ_LOW : PerformanceCounterPlugin_logic_fsm_stateNext_string = "READ_LOW ";
      PerformanceCounterPlugin_logic_fsm_CALC_LOW : PerformanceCounterPlugin_logic_fsm_stateNext_string = "CALC_LOW ";
      PerformanceCounterPlugin_logic_fsm_CSR_WRITE : PerformanceCounterPlugin_logic_fsm_stateNext_string = "CSR_WRITE";
      default : PerformanceCounterPlugin_logic_fsm_stateNext_string = "?????????";
    endcase
  end
  always @(*) begin
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_IDLE : CsrAccessPlugin_logic_fsm_stateReg_string = "IDLE      ";
      CsrAccessPlugin_logic_fsm_READ : CsrAccessPlugin_logic_fsm_stateReg_string = "READ      ";
      CsrAccessPlugin_logic_fsm_WRITE : CsrAccessPlugin_logic_fsm_stateReg_string = "WRITE     ";
      CsrAccessPlugin_logic_fsm_COMPLETION : CsrAccessPlugin_logic_fsm_stateReg_string = "COMPLETION";
      default : CsrAccessPlugin_logic_fsm_stateReg_string = "??????????";
    endcase
  end
  always @(*) begin
    case(CsrAccessPlugin_logic_fsm_stateNext)
      CsrAccessPlugin_logic_fsm_IDLE : CsrAccessPlugin_logic_fsm_stateNext_string = "IDLE      ";
      CsrAccessPlugin_logic_fsm_READ : CsrAccessPlugin_logic_fsm_stateNext_string = "READ      ";
      CsrAccessPlugin_logic_fsm_WRITE : CsrAccessPlugin_logic_fsm_stateNext_string = "WRITE     ";
      CsrAccessPlugin_logic_fsm_COMPLETION : CsrAccessPlugin_logic_fsm_stateNext_string = "COMPLETION";
      default : CsrAccessPlugin_logic_fsm_stateNext_string = "??????????";
    endcase
  end
  `endif

  always @(*) begin
    BtbPlugin_logic_ras_ptr_pop_aheadValue = BtbPlugin_logic_ras_ptr_pop;
    BtbPlugin_logic_ras_ptr_pop_aheadValue = (_zz_BtbPlugin_logic_ras_ptr_pop_aheadValue - _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_3);
  end

  assign execute_ctrl4_down_RD_ENABLE_lane0 = execute_ctrl4_RD_ENABLE_lane0_bypass;
  always @(*) begin
    execute_ctrl4_RD_ENABLE_lane0_bypass = execute_ctrl4_up_RD_ENABLE_lane0;
    if(when_ExecuteLanePlugin_l306_4) begin
      execute_ctrl4_RD_ENABLE_lane0_bypass = 1'b0;
    end
  end

  assign execute_ctrl4_down_LANE_SEL_lane0 = execute_ctrl4_LANE_SEL_lane0_bypass;
  always @(*) begin
    execute_ctrl4_LANE_SEL_lane0_bypass = execute_ctrl4_up_LANE_SEL_lane0;
    if(when_ExecuteLanePlugin_l306_4) begin
      execute_ctrl4_LANE_SEL_lane0_bypass = 1'b0;
    end
  end

  assign execute_ctrl3_down_RD_ENABLE_lane0 = execute_ctrl3_RD_ENABLE_lane0_bypass;
  always @(*) begin
    execute_ctrl3_RD_ENABLE_lane0_bypass = execute_ctrl3_up_RD_ENABLE_lane0;
    if(when_ExecuteLanePlugin_l306_3) begin
      execute_ctrl3_RD_ENABLE_lane0_bypass = 1'b0;
    end
  end

  assign execute_ctrl3_down_LANE_SEL_lane0 = execute_ctrl3_LANE_SEL_lane0_bypass;
  always @(*) begin
    execute_ctrl3_LANE_SEL_lane0_bypass = execute_ctrl3_up_LANE_SEL_lane0;
    if(when_ExecuteLanePlugin_l306_3) begin
      execute_ctrl3_LANE_SEL_lane0_bypass = 1'b0;
    end
  end

  assign execute_ctrl2_down_RD_ENABLE_lane0 = execute_ctrl2_RD_ENABLE_lane0_bypass;
  always @(*) begin
    execute_ctrl2_RD_ENABLE_lane0_bypass = execute_ctrl2_up_RD_ENABLE_lane0;
    if(when_ExecuteLanePlugin_l306_2) begin
      execute_ctrl2_RD_ENABLE_lane0_bypass = 1'b0;
    end
  end

  assign execute_ctrl2_down_LANE_SEL_lane0 = execute_ctrl2_LANE_SEL_lane0_bypass;
  always @(*) begin
    execute_ctrl2_LANE_SEL_lane0_bypass = execute_ctrl2_up_LANE_SEL_lane0;
    if(when_ExecuteLanePlugin_l306_2) begin
      execute_ctrl2_LANE_SEL_lane0_bypass = 1'b0;
    end
  end

  assign execute_ctrl1_down_RD_ENABLE_lane0 = execute_ctrl1_RD_ENABLE_lane0_bypass;
  always @(*) begin
    execute_ctrl1_RD_ENABLE_lane0_bypass = execute_ctrl1_up_RD_ENABLE_lane0;
    if(when_ExecuteLanePlugin_l306_1) begin
      execute_ctrl1_RD_ENABLE_lane0_bypass = 1'b0;
    end
  end

  assign execute_ctrl1_down_LANE_SEL_lane0 = execute_ctrl1_LANE_SEL_lane0_bypass;
  always @(*) begin
    execute_ctrl1_LANE_SEL_lane0_bypass = execute_ctrl1_up_LANE_SEL_lane0;
    if(when_ExecuteLanePlugin_l306_1) begin
      execute_ctrl1_LANE_SEL_lane0_bypass = 1'b0;
    end
  end

  assign execute_ctrl0_down_RD_ENABLE_lane0 = execute_ctrl0_RD_ENABLE_lane0_bypass;
  always @(*) begin
    execute_ctrl0_RD_ENABLE_lane0_bypass = execute_ctrl0_up_RD_ENABLE_lane0;
    if(when_ExecuteLanePlugin_l306) begin
      execute_ctrl0_RD_ENABLE_lane0_bypass = 1'b0;
    end
  end

  assign execute_ctrl0_down_LANE_SEL_lane0 = execute_ctrl0_LANE_SEL_lane0_bypass;
  always @(*) begin
    execute_ctrl0_LANE_SEL_lane0_bypass = execute_ctrl0_up_LANE_SEL_lane0;
    if(when_ExecuteLanePlugin_l306) begin
      execute_ctrl0_LANE_SEL_lane0_bypass = 1'b0;
    end
  end

  always @(*) begin
    _zz_2 = 1'b0;
    if(CsrRamPlugin_logic_writeLogic_port_valid) begin
      _zz_2 = 1'b1;
    end
  end

  always @(*) begin
    PcPlugin_logic_harts_0_aggregator_fault_1 = PcPlugin_logic_harts_0_aggregator_fault;
    if(when_PcPlugin_l80) begin
      PcPlugin_logic_harts_0_aggregator_fault_1 = _zz_PcPlugin_logic_harts_0_aggregator_fault_1_1[0];
    end
  end

  always @(*) begin
    PcPlugin_logic_harts_0_aggregator_target_1 = PcPlugin_logic_harts_0_aggregator_target;
    if(when_PcPlugin_l80) begin
      PcPlugin_logic_harts_0_aggregator_target_1 = (_zz_PcPlugin_logic_harts_0_aggregator_fault_1 ? BtbPlugin_logic_pcPort_payload_pc : 39'h0);
    end
  end

  assign decode_ctrls_1_down_LANE_SEL_0 = decode_ctrls_1_LANE_SEL_0_bypass;
  always @(*) begin
    decode_ctrls_1_LANE_SEL_0_bypass = decode_ctrls_1_up_LANE_SEL_0;
    if(decode_logic_flushes_1_onLanes_0_doIt) begin
      decode_ctrls_1_LANE_SEL_0_bypass = 1'b0;
    end
  end

  assign decode_ctrls_0_down_LANE_SEL_0 = decode_ctrls_0_LANE_SEL_0_bypass;
  always @(*) begin
    decode_ctrls_0_LANE_SEL_0_bypass = decode_ctrls_0_up_LANE_SEL_0;
    if(decode_logic_flushes_0_onLanes_0_doIt) begin
      decode_ctrls_0_LANE_SEL_0_bypass = 1'b0;
    end
  end

  assign execute_ctrl4_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 = execute_ctrl4_lane0_integer_WriteBackPlugin_logic_DATA_lane0_bypass;
  assign execute_ctrl3_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 = execute_ctrl3_lane0_integer_WriteBackPlugin_logic_DATA_lane0_bypass;
  assign execute_ctrl2_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 = execute_ctrl2_lane0_integer_WriteBackPlugin_logic_DATA_lane0_bypass;
  assign decode_ctrls_1_down_TRAP_0 = decode_ctrls_1_TRAP_0_bypass;
  always @(*) begin
    decode_ctrls_1_TRAP_0_bypass = decode_ctrls_1_up_TRAP_0;
    if(when_DecoderPlugin_l229) begin
      decode_ctrls_1_TRAP_0_bypass = 1'b1;
    end
  end

  assign execute_ctrl3_down_COMPLETED_lane0 = execute_ctrl3_COMPLETED_lane0_bypass;
  assign execute_ctrl4_down_COMPLETED_lane0 = execute_ctrl4_COMPLETED_lane0_bypass;
  assign execute_ctrl2_down_COMPLETED_lane0 = execute_ctrl2_COMPLETED_lane0_bypass;
  always @(*) begin
    early0_BranchPlugin_logic_jumpLogic_history_shifter_2 = early0_BranchPlugin_logic_jumpLogic_history_shifter_1;
    if(when_BranchPlugin_l218) begin
      early0_BranchPlugin_logic_jumpLogic_history_shifter_2 = _zz_early0_BranchPlugin_logic_jumpLogic_history_shifter_2[11 : 0];
    end
  end

  always @(*) begin
    early0_BranchPlugin_logic_jumpLogic_history_shifter_1 = early0_BranchPlugin_logic_jumpLogic_history_shifter;
    if(when_BranchPlugin_l213) begin
      early0_BranchPlugin_logic_jumpLogic_history_shifter_1 = _zz_early0_BranchPlugin_logic_jumpLogic_history_shifter_1[11 : 0];
    end
  end

  assign execute_ctrl2_down_COMMIT_lane0 = execute_ctrl2_COMMIT_lane0_bypass;
  always @(*) begin
    execute_ctrl2_COMMIT_lane0_bypass = execute_ctrl2_up_COMMIT_lane0;
    if(when_EnvPlugin_l119) begin
      if(when_EnvPlugin_l123) begin
        execute_ctrl2_COMMIT_lane0_bypass = 1'b0;
      end
    end
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_READ : begin
      end
      CsrAccessPlugin_logic_fsm_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_COMPLETION : begin
      end
      default : begin
        if(CsrAccessPlugin_logic_fsm_inject_onDecodeDo) begin
          if(CsrAccessPlugin_logic_fsm_inject_sampled) begin
            if(CsrAccessPlugin_logic_fsm_inject_trapReg) begin
              execute_ctrl2_COMMIT_lane0_bypass = 1'b0;
            end
          end
        end
      end
    endcase
  end

  assign execute_ctrl2_down_TRAP_lane0 = execute_ctrl2_TRAP_lane0_bypass;
  always @(*) begin
    execute_ctrl2_TRAP_lane0_bypass = execute_ctrl2_up_TRAP_lane0;
    if(when_EnvPlugin_l119) begin
      execute_ctrl2_TRAP_lane0_bypass = 1'b1;
    end
    if(CsrAccessPlugin_logic_fsm_inject_flushReg) begin
      execute_ctrl2_TRAP_lane0_bypass = 1'b1;
    end
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_READ : begin
      end
      CsrAccessPlugin_logic_fsm_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_COMPLETION : begin
      end
      default : begin
        if(CsrAccessPlugin_logic_fsm_inject_onDecodeDo) begin
          if(CsrAccessPlugin_logic_fsm_inject_sampled) begin
            if(CsrAccessPlugin_logic_fsm_inject_trapReg) begin
              execute_ctrl2_TRAP_lane0_bypass = 1'b1;
            end else begin
              if(CsrAccessPlugin_logic_fsm_inject_busTrapReg) begin
                execute_ctrl2_TRAP_lane0_bypass = 1'b1;
              end
            end
          end
        end
      end
    endcase
  end

  assign execute_ctrl4_down_COMMIT_lane0 = execute_ctrl4_COMMIT_lane0_bypass;
  always @(*) begin
    execute_ctrl4_COMMIT_lane0_bypass = execute_ctrl4_up_COMMIT_lane0;
    if(when_LsuPlugin_l908) begin
      if(LsuPlugin_logic_onCtrl_lsuTrap) begin
        execute_ctrl4_COMMIT_lane0_bypass = 1'b0;
      end
    end
  end

  assign execute_ctrl4_down_TRAP_lane0 = execute_ctrl4_TRAP_lane0_bypass;
  always @(*) begin
    execute_ctrl4_TRAP_lane0_bypass = execute_ctrl4_up_TRAP_lane0;
    if(when_LsuPlugin_l908) begin
      if(LsuPlugin_logic_onCtrl_lsuTrap) begin
        execute_ctrl4_TRAP_lane0_bypass = 1'b1;
      end
    end
  end

  assign execute_ctrl4_down_LsuL1_SEL_lane0 = execute_ctrl4_LsuL1_SEL_lane0_bypass;
  always @(*) begin
    execute_ctrl4_LsuL1_SEL_lane0_bypass = execute_ctrl4_up_LsuL1_SEL_lane0;
    if(when_LsuPlugin_l557_1) begin
      execute_ctrl4_LsuL1_SEL_lane0_bypass = 1'b0;
    end
  end

  assign execute_ctrl3_down_LsuL1_SEL_lane0 = execute_ctrl3_LsuL1_SEL_lane0_bypass;
  always @(*) begin
    execute_ctrl3_LsuL1_SEL_lane0_bypass = execute_ctrl3_up_LsuL1_SEL_lane0;
    if(when_LsuPlugin_l557) begin
      execute_ctrl3_LsuL1_SEL_lane0_bypass = 1'b0;
    end
  end

  assign execute_ctrl2_down_LsuPlugin_logic_FENCE_lane0 = execute_ctrl2_LsuPlugin_logic_FENCE_lane0_bypass;
  always @(*) begin
    execute_ctrl2_LsuPlugin_logic_FENCE_lane0_bypass = execute_ctrl2_up_LsuPlugin_logic_FENCE_lane0;
    if(when_LsuPlugin_l529) begin
      execute_ctrl2_LsuPlugin_logic_FENCE_lane0_bypass = 1'b0;
    end
  end

  always @(*) begin
    _zz_3 = 1'b0;
    if(BtbPlugin_logic_ras_write_valid) begin
      _zz_3 = 1'b1;
    end
  end

  always @(*) begin
    _zz_4 = 1'b0;
    if(GSharePlugin_logic_mem_writes_0_valid) begin
      _zz_4 = 1'b1;
    end
  end

  always @(*) begin
    _zz_fetch_logic_ctrls_0_haltRequest_FetchL1Plugin_l217 = 1'b0;
    if(when_FetchL1Plugin_l216) begin
      _zz_fetch_logic_ctrls_0_haltRequest_FetchL1Plugin_l217 = 1'b1;
    end
  end

  always @(*) begin
    _zz_5 = 1'b0;
    if(FetchL1Plugin_logic_plru_write_valid) begin
      _zz_5 = 1'b1;
    end
  end

  always @(*) begin
    _zz_6 = 1'b0;
    if(FetchL1Plugin_logic_banks_1_write_valid) begin
      _zz_6 = 1'b1;
    end
  end

  always @(*) begin
    _zz_7 = 1'b0;
    if(FetchL1Plugin_logic_banks_0_write_valid) begin
      _zz_7 = 1'b1;
    end
  end

  assign execute_ctrl3_down_LsuL1Plugin_logic_SHARED_lane0_plru_0 = execute_ctrl3_LsuL1Plugin_logic_SHARED_lane0_bypass_plru_0;
  assign execute_ctrl3_down_LsuL1Plugin_logic_SHARED_lane0_dirty = execute_ctrl3_LsuL1Plugin_logic_SHARED_lane0_bypass_dirty;
  assign execute_ctrl4_down_LsuL1Plugin_logic_FREEZE_HAZARD_lane0 = execute_ctrl4_LsuL1Plugin_logic_FREEZE_HAZARD_lane0_bypass;
  assign execute_ctrl3_down_LsuL1Plugin_logic_FREEZE_HAZARD_lane0 = execute_ctrl3_LsuL1Plugin_logic_FREEZE_HAZARD_lane0_bypass;
  always @(*) begin
    _zz_8 = 1'b0;
    if(LsuL1Plugin_logic_writeback_read_slotReadLast_valid) begin
      _zz_8 = 1'b1;
    end
  end

  always @(*) begin
    _zz_9 = 1'b0;
    if(LsuL1Plugin_logic_shared_write_valid) begin
      _zz_9 = 1'b1;
    end
  end

  assign AlignerPlugin_api_singleFetch = 1'b0;
  assign AlignerPlugin_api_haltIt = 1'b0;
  always @(*) begin
    DispatchPlugin_api_haltDispatch = 1'b0;
    if(LsuPlugin_logic_onAddress0_access_sbWaiter) begin
      DispatchPlugin_api_haltDispatch = 1'b1;
    end
    if(LsuPlugin_logic_onCtrl_hartRegulation_valid) begin
      DispatchPlugin_api_haltDispatch = 1'b1;
    end
  end

  always @(*) begin
    CsrRamPlugin_api_holdRead = 1'b0;
    if(PerformanceCounterPlugin_logic_csrRead_requested) begin
      if(when_PerformanceCounterPlugin_l342) begin
        CsrRamPlugin_api_holdRead = 1'b1;
      end
    end
  end

  always @(*) begin
    CsrRamPlugin_api_holdWrite = 1'b0;
    if(PerformanceCounterPlugin_logic_fsm_holdCsrWrite) begin
      CsrRamPlugin_api_holdWrite = 1'b1;
    end
  end

  always @(*) begin
    TrapPlugin_api_harts_0_redo = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
        if(!when_TrapPlugin_l453) begin
          case(TrapPlugin_logic_harts_0_trap_pending_state_code)
            4'b0000 : begin
            end
            4'b0001 : begin
            end
            4'b0010 : begin
            end
            4'b0100 : begin
              TrapPlugin_api_harts_0_redo = 1'b1;
            end
            4'b0101 : begin
            end
            4'b1000 : begin
            end
            4'b0110 : begin
            end
            4'b0111 : begin
            end
            default : begin
            end
          endcase
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_WAIT : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
        if(TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_valid) begin
          TrapPlugin_api_harts_0_redo = 1'b1;
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_api_harts_0_askWake = 1'b0;
    if(when_TrapPlugin_l269) begin
      TrapPlugin_api_harts_0_askWake = 1'b1;
    end
  end

  always @(*) begin
    TrapPlugin_api_harts_0_rvTrap = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_WAIT : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
        TrapPlugin_api_harts_0_rvTrap = 1'b1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  assign TrapPlugin_api_harts_0_holdPrivChange = 1'b0;
  always @(*) begin
    PmpPlugin_logic_entries_0_cfgNext_kind = PmpPlugin_logic_entries_0_cfg_kind;
    if(when_CsrAccessPlugin_l352_4) begin
      PmpPlugin_logic_entries_0_cfgNext_kind = CsrAccessPlugin_bus_write_bits[4 : 3];
    end
  end

  always @(*) begin
    PmpPlugin_logic_entries_0_cfgNext_read = PmpPlugin_logic_entries_0_cfg_read;
    if(when_CsrAccessPlugin_l352_4) begin
      PmpPlugin_logic_entries_0_cfgNext_read = CsrAccessPlugin_bus_write_bits[0];
    end
  end

  always @(*) begin
    PmpPlugin_logic_entries_0_cfgNext_write = PmpPlugin_logic_entries_0_cfg_write;
    if(when_CsrAccessPlugin_l352_4) begin
      PmpPlugin_logic_entries_0_cfgNext_write = CsrAccessPlugin_bus_write_bits[1];
    end
  end

  always @(*) begin
    PmpPlugin_logic_entries_0_cfgNext_execute = PmpPlugin_logic_entries_0_cfg_execute;
    if(when_CsrAccessPlugin_l352_4) begin
      PmpPlugin_logic_entries_0_cfgNext_execute = CsrAccessPlugin_bus_write_bits[2];
    end
  end

  always @(*) begin
    PmpPlugin_logic_entries_0_cfgNext_locked = PmpPlugin_logic_entries_0_cfg_locked;
    if(when_CsrAccessPlugin_l352_4) begin
      PmpPlugin_logic_entries_0_cfgNext_locked = CsrAccessPlugin_bus_write_bits[7];
    end
  end

  assign when_PmpPlugin_l127 = (! PmpPlugin_logic_entries_0_cfg_locked);
  assign when_PmpPlugin_l129 = (! PmpPlugin_logic_entries_0_cfgNext_read);
  assign _zz_PmpPlugin_logic_entries_0_napot = (~ PmpPlugin_logic_entries_0_address[19 : 0]);
  assign _zz_PmpPlugin_logic_entries_0_napot_1 = _zz_PmpPlugin_logic_entries_0_napot[0];
  assign _zz_PmpPlugin_logic_entries_0_napot_2 = _zz_PmpPlugin_logic_entries_0_napot[1];
  assign _zz_PmpPlugin_logic_entries_0_napot_3 = _zz_PmpPlugin_logic_entries_0_napot[2];
  assign _zz_PmpPlugin_logic_entries_0_napot_4 = _zz_PmpPlugin_logic_entries_0_napot[4];
  assign _zz_PmpPlugin_logic_entries_0_napot_5 = _zz_PmpPlugin_logic_entries_0_napot[5];
  assign _zz_PmpPlugin_logic_entries_0_napot_6 = _zz_PmpPlugin_logic_entries_0_napot[6];
  assign _zz_PmpPlugin_logic_entries_0_napot_7 = _zz_PmpPlugin_logic_entries_0_napot[8];
  assign _zz_PmpPlugin_logic_entries_0_napot_8 = _zz_PmpPlugin_logic_entries_0_napot[9];
  assign _zz_PmpPlugin_logic_entries_0_napot_9 = _zz_PmpPlugin_logic_entries_0_napot[10];
  assign _zz_PmpPlugin_logic_entries_0_napot_10 = _zz_PmpPlugin_logic_entries_0_napot[12];
  assign _zz_PmpPlugin_logic_entries_0_napot_11 = _zz_PmpPlugin_logic_entries_0_napot[13];
  assign _zz_PmpPlugin_logic_entries_0_napot_12 = _zz_PmpPlugin_logic_entries_0_napot[14];
  assign _zz_PmpPlugin_logic_entries_0_napot_13 = _zz_PmpPlugin_logic_entries_0_napot[16];
  assign _zz_PmpPlugin_logic_entries_0_napot_14 = _zz_PmpPlugin_logic_entries_0_napot[17];
  assign _zz_PmpPlugin_logic_entries_0_napot_15 = _zz_PmpPlugin_logic_entries_0_napot[18];
  always @(*) begin
    _zz_PmpPlugin_logic_entries_0_napot_16[0] = _zz_PmpPlugin_logic_entries_0_napot_1;
    _zz_PmpPlugin_logic_entries_0_napot_16[1] = (|{_zz_PmpPlugin_logic_entries_0_napot_2,_zz_PmpPlugin_logic_entries_0_napot_1});
    _zz_PmpPlugin_logic_entries_0_napot_16[2] = (|{_zz_PmpPlugin_logic_entries_0_napot_3,{_zz_PmpPlugin_logic_entries_0_napot_2,_zz_PmpPlugin_logic_entries_0_napot_1}});
    _zz_PmpPlugin_logic_entries_0_napot_16[3] = _zz_PmpPlugin_logic_entries_0_napot_17;
    _zz_PmpPlugin_logic_entries_0_napot_16[4] = (_zz_PmpPlugin_logic_entries_0_napot_4 || _zz_PmpPlugin_logic_entries_0_napot_17);
    _zz_PmpPlugin_logic_entries_0_napot_16[5] = ((|{_zz_PmpPlugin_logic_entries_0_napot_5,_zz_PmpPlugin_logic_entries_0_napot_4}) || _zz_PmpPlugin_logic_entries_0_napot_17);
    _zz_PmpPlugin_logic_entries_0_napot_16[6] = ((|{_zz_PmpPlugin_logic_entries_0_napot_6,{_zz_PmpPlugin_logic_entries_0_napot_5,_zz_PmpPlugin_logic_entries_0_napot_4}}) || _zz_PmpPlugin_logic_entries_0_napot_17);
    _zz_PmpPlugin_logic_entries_0_napot_16[7] = (_zz_PmpPlugin_logic_entries_0_napot_18 || _zz_PmpPlugin_logic_entries_0_napot_17);
    _zz_PmpPlugin_logic_entries_0_napot_16[8] = (_zz_PmpPlugin_logic_entries_0_napot_7 || _zz_PmpPlugin_logic_entries_0_napot_19);
    _zz_PmpPlugin_logic_entries_0_napot_16[9] = ((|{_zz_PmpPlugin_logic_entries_0_napot_8,_zz_PmpPlugin_logic_entries_0_napot_7}) || _zz_PmpPlugin_logic_entries_0_napot_19);
    _zz_PmpPlugin_logic_entries_0_napot_16[10] = ((|{_zz_PmpPlugin_logic_entries_0_napot_9,{_zz_PmpPlugin_logic_entries_0_napot_8,_zz_PmpPlugin_logic_entries_0_napot_7}}) || _zz_PmpPlugin_logic_entries_0_napot_19);
    _zz_PmpPlugin_logic_entries_0_napot_16[11] = (_zz_PmpPlugin_logic_entries_0_napot_20 || _zz_PmpPlugin_logic_entries_0_napot_19);
    _zz_PmpPlugin_logic_entries_0_napot_16[12] = (_zz_PmpPlugin_logic_entries_0_napot_10 || _zz_PmpPlugin_logic_entries_0_napot_21);
    _zz_PmpPlugin_logic_entries_0_napot_16[13] = ((|{_zz_PmpPlugin_logic_entries_0_napot_11,_zz_PmpPlugin_logic_entries_0_napot_10}) || _zz_PmpPlugin_logic_entries_0_napot_21);
    _zz_PmpPlugin_logic_entries_0_napot_16[14] = ((|{_zz_PmpPlugin_logic_entries_0_napot_12,{_zz_PmpPlugin_logic_entries_0_napot_11,_zz_PmpPlugin_logic_entries_0_napot_10}}) || _zz_PmpPlugin_logic_entries_0_napot_21);
    _zz_PmpPlugin_logic_entries_0_napot_16[15] = (_zz_PmpPlugin_logic_entries_0_napot_22 || _zz_PmpPlugin_logic_entries_0_napot_21);
    _zz_PmpPlugin_logic_entries_0_napot_16[16] = (_zz_PmpPlugin_logic_entries_0_napot_13 || _zz_PmpPlugin_logic_entries_0_napot_23);
    _zz_PmpPlugin_logic_entries_0_napot_16[17] = ((|{_zz_PmpPlugin_logic_entries_0_napot_14,_zz_PmpPlugin_logic_entries_0_napot_13}) || _zz_PmpPlugin_logic_entries_0_napot_23);
    _zz_PmpPlugin_logic_entries_0_napot_16[18] = ((|{_zz_PmpPlugin_logic_entries_0_napot_15,{_zz_PmpPlugin_logic_entries_0_napot_14,_zz_PmpPlugin_logic_entries_0_napot_13}}) || _zz_PmpPlugin_logic_entries_0_napot_23);
    _zz_PmpPlugin_logic_entries_0_napot_16[19] = ((|{_zz_PmpPlugin_logic_entries_0_napot[19],{_zz_PmpPlugin_logic_entries_0_napot_15,{_zz_PmpPlugin_logic_entries_0_napot_14,_zz_PmpPlugin_logic_entries_0_napot_13}}}) || _zz_PmpPlugin_logic_entries_0_napot_23);
  end

  assign _zz_PmpPlugin_logic_entries_0_napot_17 = (|{_zz_PmpPlugin_logic_entries_0_napot[3],{_zz_PmpPlugin_logic_entries_0_napot_3,{_zz_PmpPlugin_logic_entries_0_napot_2,_zz_PmpPlugin_logic_entries_0_napot_1}}});
  assign _zz_PmpPlugin_logic_entries_0_napot_18 = (|{_zz_PmpPlugin_logic_entries_0_napot[7],{_zz_PmpPlugin_logic_entries_0_napot_6,{_zz_PmpPlugin_logic_entries_0_napot_5,_zz_PmpPlugin_logic_entries_0_napot_4}}});
  assign _zz_PmpPlugin_logic_entries_0_napot_19 = (|{_zz_PmpPlugin_logic_entries_0_napot_18,_zz_PmpPlugin_logic_entries_0_napot_17});
  assign _zz_PmpPlugin_logic_entries_0_napot_20 = (|{_zz_PmpPlugin_logic_entries_0_napot[11],{_zz_PmpPlugin_logic_entries_0_napot_9,{_zz_PmpPlugin_logic_entries_0_napot_8,_zz_PmpPlugin_logic_entries_0_napot_7}}});
  assign _zz_PmpPlugin_logic_entries_0_napot_21 = (|{_zz_PmpPlugin_logic_entries_0_napot_20,{_zz_PmpPlugin_logic_entries_0_napot_18,_zz_PmpPlugin_logic_entries_0_napot_17}});
  assign _zz_PmpPlugin_logic_entries_0_napot_22 = (|{_zz_PmpPlugin_logic_entries_0_napot[15],{_zz_PmpPlugin_logic_entries_0_napot_12,{_zz_PmpPlugin_logic_entries_0_napot_11,_zz_PmpPlugin_logic_entries_0_napot_10}}});
  assign _zz_PmpPlugin_logic_entries_0_napot_23 = (|{_zz_PmpPlugin_logic_entries_0_napot_22,{_zz_PmpPlugin_logic_entries_0_napot_20,{_zz_PmpPlugin_logic_entries_0_napot_18,_zz_PmpPlugin_logic_entries_0_napot_17}}});
  assign PmpPlugin_logic_entries_0_napot = _zz_PmpPlugin_logic_entries_0_napot_24[20 : 1];
  always @(*) begin
    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4 = (PmpPlugin_logic_entries_0_isNapot ? 10'h3ff : 10'h0);
    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4[9] = (PmpPlugin_logic_entries_0_address[0] && PmpPlugin_logic_entries_0_isNapot);
  end

  always @(*) begin
    PmpPlugin_logic_entries_1_cfgNext_kind = PmpPlugin_logic_entries_1_cfg_kind;
    if(when_CsrAccessPlugin_l352_4) begin
      PmpPlugin_logic_entries_1_cfgNext_kind = CsrAccessPlugin_bus_write_bits[12 : 11];
    end
  end

  always @(*) begin
    PmpPlugin_logic_entries_1_cfgNext_read = PmpPlugin_logic_entries_1_cfg_read;
    if(when_CsrAccessPlugin_l352_4) begin
      PmpPlugin_logic_entries_1_cfgNext_read = CsrAccessPlugin_bus_write_bits[8];
    end
  end

  always @(*) begin
    PmpPlugin_logic_entries_1_cfgNext_write = PmpPlugin_logic_entries_1_cfg_write;
    if(when_CsrAccessPlugin_l352_4) begin
      PmpPlugin_logic_entries_1_cfgNext_write = CsrAccessPlugin_bus_write_bits[9];
    end
  end

  always @(*) begin
    PmpPlugin_logic_entries_1_cfgNext_execute = PmpPlugin_logic_entries_1_cfg_execute;
    if(when_CsrAccessPlugin_l352_4) begin
      PmpPlugin_logic_entries_1_cfgNext_execute = CsrAccessPlugin_bus_write_bits[10];
    end
  end

  always @(*) begin
    PmpPlugin_logic_entries_1_cfgNext_locked = PmpPlugin_logic_entries_1_cfg_locked;
    if(when_CsrAccessPlugin_l352_4) begin
      PmpPlugin_logic_entries_1_cfgNext_locked = CsrAccessPlugin_bus_write_bits[15];
    end
  end

  assign when_PmpPlugin_l127_1 = (! PmpPlugin_logic_entries_1_cfg_locked);
  assign when_PmpPlugin_l129_1 = (! PmpPlugin_logic_entries_1_cfgNext_read);
  assign _zz_PmpPlugin_logic_entries_1_napot = (~ PmpPlugin_logic_entries_1_address[19 : 0]);
  assign _zz_PmpPlugin_logic_entries_1_napot_1 = _zz_PmpPlugin_logic_entries_1_napot[0];
  assign _zz_PmpPlugin_logic_entries_1_napot_2 = _zz_PmpPlugin_logic_entries_1_napot[1];
  assign _zz_PmpPlugin_logic_entries_1_napot_3 = _zz_PmpPlugin_logic_entries_1_napot[2];
  assign _zz_PmpPlugin_logic_entries_1_napot_4 = _zz_PmpPlugin_logic_entries_1_napot[4];
  assign _zz_PmpPlugin_logic_entries_1_napot_5 = _zz_PmpPlugin_logic_entries_1_napot[5];
  assign _zz_PmpPlugin_logic_entries_1_napot_6 = _zz_PmpPlugin_logic_entries_1_napot[6];
  assign _zz_PmpPlugin_logic_entries_1_napot_7 = _zz_PmpPlugin_logic_entries_1_napot[8];
  assign _zz_PmpPlugin_logic_entries_1_napot_8 = _zz_PmpPlugin_logic_entries_1_napot[9];
  assign _zz_PmpPlugin_logic_entries_1_napot_9 = _zz_PmpPlugin_logic_entries_1_napot[10];
  assign _zz_PmpPlugin_logic_entries_1_napot_10 = _zz_PmpPlugin_logic_entries_1_napot[12];
  assign _zz_PmpPlugin_logic_entries_1_napot_11 = _zz_PmpPlugin_logic_entries_1_napot[13];
  assign _zz_PmpPlugin_logic_entries_1_napot_12 = _zz_PmpPlugin_logic_entries_1_napot[14];
  assign _zz_PmpPlugin_logic_entries_1_napot_13 = _zz_PmpPlugin_logic_entries_1_napot[16];
  assign _zz_PmpPlugin_logic_entries_1_napot_14 = _zz_PmpPlugin_logic_entries_1_napot[17];
  assign _zz_PmpPlugin_logic_entries_1_napot_15 = _zz_PmpPlugin_logic_entries_1_napot[18];
  always @(*) begin
    _zz_PmpPlugin_logic_entries_1_napot_16[0] = _zz_PmpPlugin_logic_entries_1_napot_1;
    _zz_PmpPlugin_logic_entries_1_napot_16[1] = (|{_zz_PmpPlugin_logic_entries_1_napot_2,_zz_PmpPlugin_logic_entries_1_napot_1});
    _zz_PmpPlugin_logic_entries_1_napot_16[2] = (|{_zz_PmpPlugin_logic_entries_1_napot_3,{_zz_PmpPlugin_logic_entries_1_napot_2,_zz_PmpPlugin_logic_entries_1_napot_1}});
    _zz_PmpPlugin_logic_entries_1_napot_16[3] = _zz_PmpPlugin_logic_entries_1_napot_17;
    _zz_PmpPlugin_logic_entries_1_napot_16[4] = (_zz_PmpPlugin_logic_entries_1_napot_4 || _zz_PmpPlugin_logic_entries_1_napot_17);
    _zz_PmpPlugin_logic_entries_1_napot_16[5] = ((|{_zz_PmpPlugin_logic_entries_1_napot_5,_zz_PmpPlugin_logic_entries_1_napot_4}) || _zz_PmpPlugin_logic_entries_1_napot_17);
    _zz_PmpPlugin_logic_entries_1_napot_16[6] = ((|{_zz_PmpPlugin_logic_entries_1_napot_6,{_zz_PmpPlugin_logic_entries_1_napot_5,_zz_PmpPlugin_logic_entries_1_napot_4}}) || _zz_PmpPlugin_logic_entries_1_napot_17);
    _zz_PmpPlugin_logic_entries_1_napot_16[7] = (_zz_PmpPlugin_logic_entries_1_napot_18 || _zz_PmpPlugin_logic_entries_1_napot_17);
    _zz_PmpPlugin_logic_entries_1_napot_16[8] = (_zz_PmpPlugin_logic_entries_1_napot_7 || _zz_PmpPlugin_logic_entries_1_napot_19);
    _zz_PmpPlugin_logic_entries_1_napot_16[9] = ((|{_zz_PmpPlugin_logic_entries_1_napot_8,_zz_PmpPlugin_logic_entries_1_napot_7}) || _zz_PmpPlugin_logic_entries_1_napot_19);
    _zz_PmpPlugin_logic_entries_1_napot_16[10] = ((|{_zz_PmpPlugin_logic_entries_1_napot_9,{_zz_PmpPlugin_logic_entries_1_napot_8,_zz_PmpPlugin_logic_entries_1_napot_7}}) || _zz_PmpPlugin_logic_entries_1_napot_19);
    _zz_PmpPlugin_logic_entries_1_napot_16[11] = (_zz_PmpPlugin_logic_entries_1_napot_20 || _zz_PmpPlugin_logic_entries_1_napot_19);
    _zz_PmpPlugin_logic_entries_1_napot_16[12] = (_zz_PmpPlugin_logic_entries_1_napot_10 || _zz_PmpPlugin_logic_entries_1_napot_21);
    _zz_PmpPlugin_logic_entries_1_napot_16[13] = ((|{_zz_PmpPlugin_logic_entries_1_napot_11,_zz_PmpPlugin_logic_entries_1_napot_10}) || _zz_PmpPlugin_logic_entries_1_napot_21);
    _zz_PmpPlugin_logic_entries_1_napot_16[14] = ((|{_zz_PmpPlugin_logic_entries_1_napot_12,{_zz_PmpPlugin_logic_entries_1_napot_11,_zz_PmpPlugin_logic_entries_1_napot_10}}) || _zz_PmpPlugin_logic_entries_1_napot_21);
    _zz_PmpPlugin_logic_entries_1_napot_16[15] = (_zz_PmpPlugin_logic_entries_1_napot_22 || _zz_PmpPlugin_logic_entries_1_napot_21);
    _zz_PmpPlugin_logic_entries_1_napot_16[16] = (_zz_PmpPlugin_logic_entries_1_napot_13 || _zz_PmpPlugin_logic_entries_1_napot_23);
    _zz_PmpPlugin_logic_entries_1_napot_16[17] = ((|{_zz_PmpPlugin_logic_entries_1_napot_14,_zz_PmpPlugin_logic_entries_1_napot_13}) || _zz_PmpPlugin_logic_entries_1_napot_23);
    _zz_PmpPlugin_logic_entries_1_napot_16[18] = ((|{_zz_PmpPlugin_logic_entries_1_napot_15,{_zz_PmpPlugin_logic_entries_1_napot_14,_zz_PmpPlugin_logic_entries_1_napot_13}}) || _zz_PmpPlugin_logic_entries_1_napot_23);
    _zz_PmpPlugin_logic_entries_1_napot_16[19] = ((|{_zz_PmpPlugin_logic_entries_1_napot[19],{_zz_PmpPlugin_logic_entries_1_napot_15,{_zz_PmpPlugin_logic_entries_1_napot_14,_zz_PmpPlugin_logic_entries_1_napot_13}}}) || _zz_PmpPlugin_logic_entries_1_napot_23);
  end

  assign _zz_PmpPlugin_logic_entries_1_napot_17 = (|{_zz_PmpPlugin_logic_entries_1_napot[3],{_zz_PmpPlugin_logic_entries_1_napot_3,{_zz_PmpPlugin_logic_entries_1_napot_2,_zz_PmpPlugin_logic_entries_1_napot_1}}});
  assign _zz_PmpPlugin_logic_entries_1_napot_18 = (|{_zz_PmpPlugin_logic_entries_1_napot[7],{_zz_PmpPlugin_logic_entries_1_napot_6,{_zz_PmpPlugin_logic_entries_1_napot_5,_zz_PmpPlugin_logic_entries_1_napot_4}}});
  assign _zz_PmpPlugin_logic_entries_1_napot_19 = (|{_zz_PmpPlugin_logic_entries_1_napot_18,_zz_PmpPlugin_logic_entries_1_napot_17});
  assign _zz_PmpPlugin_logic_entries_1_napot_20 = (|{_zz_PmpPlugin_logic_entries_1_napot[11],{_zz_PmpPlugin_logic_entries_1_napot_9,{_zz_PmpPlugin_logic_entries_1_napot_8,_zz_PmpPlugin_logic_entries_1_napot_7}}});
  assign _zz_PmpPlugin_logic_entries_1_napot_21 = (|{_zz_PmpPlugin_logic_entries_1_napot_20,{_zz_PmpPlugin_logic_entries_1_napot_18,_zz_PmpPlugin_logic_entries_1_napot_17}});
  assign _zz_PmpPlugin_logic_entries_1_napot_22 = (|{_zz_PmpPlugin_logic_entries_1_napot[15],{_zz_PmpPlugin_logic_entries_1_napot_12,{_zz_PmpPlugin_logic_entries_1_napot_11,_zz_PmpPlugin_logic_entries_1_napot_10}}});
  assign _zz_PmpPlugin_logic_entries_1_napot_23 = (|{_zz_PmpPlugin_logic_entries_1_napot_22,{_zz_PmpPlugin_logic_entries_1_napot_20,{_zz_PmpPlugin_logic_entries_1_napot_18,_zz_PmpPlugin_logic_entries_1_napot_17}}});
  assign PmpPlugin_logic_entries_1_napot = _zz_PmpPlugin_logic_entries_1_napot_24[20 : 1];
  always @(*) begin
    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_7 = (PmpPlugin_logic_entries_1_isNapot ? 10'h3ff : 10'h0);
    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_7[9] = (PmpPlugin_logic_entries_1_address[0] && PmpPlugin_logic_entries_1_isNapot);
  end

  always @(*) begin
    PmpPlugin_logic_entries_2_cfgNext_kind = PmpPlugin_logic_entries_2_cfg_kind;
    if(when_CsrAccessPlugin_l352_4) begin
      PmpPlugin_logic_entries_2_cfgNext_kind = CsrAccessPlugin_bus_write_bits[20 : 19];
    end
  end

  always @(*) begin
    PmpPlugin_logic_entries_2_cfgNext_read = PmpPlugin_logic_entries_2_cfg_read;
    if(when_CsrAccessPlugin_l352_4) begin
      PmpPlugin_logic_entries_2_cfgNext_read = CsrAccessPlugin_bus_write_bits[16];
    end
  end

  always @(*) begin
    PmpPlugin_logic_entries_2_cfgNext_write = PmpPlugin_logic_entries_2_cfg_write;
    if(when_CsrAccessPlugin_l352_4) begin
      PmpPlugin_logic_entries_2_cfgNext_write = CsrAccessPlugin_bus_write_bits[17];
    end
  end

  always @(*) begin
    PmpPlugin_logic_entries_2_cfgNext_execute = PmpPlugin_logic_entries_2_cfg_execute;
    if(when_CsrAccessPlugin_l352_4) begin
      PmpPlugin_logic_entries_2_cfgNext_execute = CsrAccessPlugin_bus_write_bits[18];
    end
  end

  always @(*) begin
    PmpPlugin_logic_entries_2_cfgNext_locked = PmpPlugin_logic_entries_2_cfg_locked;
    if(when_CsrAccessPlugin_l352_4) begin
      PmpPlugin_logic_entries_2_cfgNext_locked = CsrAccessPlugin_bus_write_bits[23];
    end
  end

  assign when_PmpPlugin_l127_2 = (! PmpPlugin_logic_entries_2_cfg_locked);
  assign when_PmpPlugin_l129_2 = (! PmpPlugin_logic_entries_2_cfgNext_read);
  assign _zz_PmpPlugin_logic_entries_2_napot = (~ PmpPlugin_logic_entries_2_address[19 : 0]);
  assign _zz_PmpPlugin_logic_entries_2_napot_1 = _zz_PmpPlugin_logic_entries_2_napot[0];
  assign _zz_PmpPlugin_logic_entries_2_napot_2 = _zz_PmpPlugin_logic_entries_2_napot[1];
  assign _zz_PmpPlugin_logic_entries_2_napot_3 = _zz_PmpPlugin_logic_entries_2_napot[2];
  assign _zz_PmpPlugin_logic_entries_2_napot_4 = _zz_PmpPlugin_logic_entries_2_napot[4];
  assign _zz_PmpPlugin_logic_entries_2_napot_5 = _zz_PmpPlugin_logic_entries_2_napot[5];
  assign _zz_PmpPlugin_logic_entries_2_napot_6 = _zz_PmpPlugin_logic_entries_2_napot[6];
  assign _zz_PmpPlugin_logic_entries_2_napot_7 = _zz_PmpPlugin_logic_entries_2_napot[8];
  assign _zz_PmpPlugin_logic_entries_2_napot_8 = _zz_PmpPlugin_logic_entries_2_napot[9];
  assign _zz_PmpPlugin_logic_entries_2_napot_9 = _zz_PmpPlugin_logic_entries_2_napot[10];
  assign _zz_PmpPlugin_logic_entries_2_napot_10 = _zz_PmpPlugin_logic_entries_2_napot[12];
  assign _zz_PmpPlugin_logic_entries_2_napot_11 = _zz_PmpPlugin_logic_entries_2_napot[13];
  assign _zz_PmpPlugin_logic_entries_2_napot_12 = _zz_PmpPlugin_logic_entries_2_napot[14];
  assign _zz_PmpPlugin_logic_entries_2_napot_13 = _zz_PmpPlugin_logic_entries_2_napot[16];
  assign _zz_PmpPlugin_logic_entries_2_napot_14 = _zz_PmpPlugin_logic_entries_2_napot[17];
  assign _zz_PmpPlugin_logic_entries_2_napot_15 = _zz_PmpPlugin_logic_entries_2_napot[18];
  always @(*) begin
    _zz_PmpPlugin_logic_entries_2_napot_16[0] = _zz_PmpPlugin_logic_entries_2_napot_1;
    _zz_PmpPlugin_logic_entries_2_napot_16[1] = (|{_zz_PmpPlugin_logic_entries_2_napot_2,_zz_PmpPlugin_logic_entries_2_napot_1});
    _zz_PmpPlugin_logic_entries_2_napot_16[2] = (|{_zz_PmpPlugin_logic_entries_2_napot_3,{_zz_PmpPlugin_logic_entries_2_napot_2,_zz_PmpPlugin_logic_entries_2_napot_1}});
    _zz_PmpPlugin_logic_entries_2_napot_16[3] = _zz_PmpPlugin_logic_entries_2_napot_17;
    _zz_PmpPlugin_logic_entries_2_napot_16[4] = (_zz_PmpPlugin_logic_entries_2_napot_4 || _zz_PmpPlugin_logic_entries_2_napot_17);
    _zz_PmpPlugin_logic_entries_2_napot_16[5] = ((|{_zz_PmpPlugin_logic_entries_2_napot_5,_zz_PmpPlugin_logic_entries_2_napot_4}) || _zz_PmpPlugin_logic_entries_2_napot_17);
    _zz_PmpPlugin_logic_entries_2_napot_16[6] = ((|{_zz_PmpPlugin_logic_entries_2_napot_6,{_zz_PmpPlugin_logic_entries_2_napot_5,_zz_PmpPlugin_logic_entries_2_napot_4}}) || _zz_PmpPlugin_logic_entries_2_napot_17);
    _zz_PmpPlugin_logic_entries_2_napot_16[7] = (_zz_PmpPlugin_logic_entries_2_napot_18 || _zz_PmpPlugin_logic_entries_2_napot_17);
    _zz_PmpPlugin_logic_entries_2_napot_16[8] = (_zz_PmpPlugin_logic_entries_2_napot_7 || _zz_PmpPlugin_logic_entries_2_napot_19);
    _zz_PmpPlugin_logic_entries_2_napot_16[9] = ((|{_zz_PmpPlugin_logic_entries_2_napot_8,_zz_PmpPlugin_logic_entries_2_napot_7}) || _zz_PmpPlugin_logic_entries_2_napot_19);
    _zz_PmpPlugin_logic_entries_2_napot_16[10] = ((|{_zz_PmpPlugin_logic_entries_2_napot_9,{_zz_PmpPlugin_logic_entries_2_napot_8,_zz_PmpPlugin_logic_entries_2_napot_7}}) || _zz_PmpPlugin_logic_entries_2_napot_19);
    _zz_PmpPlugin_logic_entries_2_napot_16[11] = (_zz_PmpPlugin_logic_entries_2_napot_20 || _zz_PmpPlugin_logic_entries_2_napot_19);
    _zz_PmpPlugin_logic_entries_2_napot_16[12] = (_zz_PmpPlugin_logic_entries_2_napot_10 || _zz_PmpPlugin_logic_entries_2_napot_21);
    _zz_PmpPlugin_logic_entries_2_napot_16[13] = ((|{_zz_PmpPlugin_logic_entries_2_napot_11,_zz_PmpPlugin_logic_entries_2_napot_10}) || _zz_PmpPlugin_logic_entries_2_napot_21);
    _zz_PmpPlugin_logic_entries_2_napot_16[14] = ((|{_zz_PmpPlugin_logic_entries_2_napot_12,{_zz_PmpPlugin_logic_entries_2_napot_11,_zz_PmpPlugin_logic_entries_2_napot_10}}) || _zz_PmpPlugin_logic_entries_2_napot_21);
    _zz_PmpPlugin_logic_entries_2_napot_16[15] = (_zz_PmpPlugin_logic_entries_2_napot_22 || _zz_PmpPlugin_logic_entries_2_napot_21);
    _zz_PmpPlugin_logic_entries_2_napot_16[16] = (_zz_PmpPlugin_logic_entries_2_napot_13 || _zz_PmpPlugin_logic_entries_2_napot_23);
    _zz_PmpPlugin_logic_entries_2_napot_16[17] = ((|{_zz_PmpPlugin_logic_entries_2_napot_14,_zz_PmpPlugin_logic_entries_2_napot_13}) || _zz_PmpPlugin_logic_entries_2_napot_23);
    _zz_PmpPlugin_logic_entries_2_napot_16[18] = ((|{_zz_PmpPlugin_logic_entries_2_napot_15,{_zz_PmpPlugin_logic_entries_2_napot_14,_zz_PmpPlugin_logic_entries_2_napot_13}}) || _zz_PmpPlugin_logic_entries_2_napot_23);
    _zz_PmpPlugin_logic_entries_2_napot_16[19] = ((|{_zz_PmpPlugin_logic_entries_2_napot[19],{_zz_PmpPlugin_logic_entries_2_napot_15,{_zz_PmpPlugin_logic_entries_2_napot_14,_zz_PmpPlugin_logic_entries_2_napot_13}}}) || _zz_PmpPlugin_logic_entries_2_napot_23);
  end

  assign _zz_PmpPlugin_logic_entries_2_napot_17 = (|{_zz_PmpPlugin_logic_entries_2_napot[3],{_zz_PmpPlugin_logic_entries_2_napot_3,{_zz_PmpPlugin_logic_entries_2_napot_2,_zz_PmpPlugin_logic_entries_2_napot_1}}});
  assign _zz_PmpPlugin_logic_entries_2_napot_18 = (|{_zz_PmpPlugin_logic_entries_2_napot[7],{_zz_PmpPlugin_logic_entries_2_napot_6,{_zz_PmpPlugin_logic_entries_2_napot_5,_zz_PmpPlugin_logic_entries_2_napot_4}}});
  assign _zz_PmpPlugin_logic_entries_2_napot_19 = (|{_zz_PmpPlugin_logic_entries_2_napot_18,_zz_PmpPlugin_logic_entries_2_napot_17});
  assign _zz_PmpPlugin_logic_entries_2_napot_20 = (|{_zz_PmpPlugin_logic_entries_2_napot[11],{_zz_PmpPlugin_logic_entries_2_napot_9,{_zz_PmpPlugin_logic_entries_2_napot_8,_zz_PmpPlugin_logic_entries_2_napot_7}}});
  assign _zz_PmpPlugin_logic_entries_2_napot_21 = (|{_zz_PmpPlugin_logic_entries_2_napot_20,{_zz_PmpPlugin_logic_entries_2_napot_18,_zz_PmpPlugin_logic_entries_2_napot_17}});
  assign _zz_PmpPlugin_logic_entries_2_napot_22 = (|{_zz_PmpPlugin_logic_entries_2_napot[15],{_zz_PmpPlugin_logic_entries_2_napot_12,{_zz_PmpPlugin_logic_entries_2_napot_11,_zz_PmpPlugin_logic_entries_2_napot_10}}});
  assign _zz_PmpPlugin_logic_entries_2_napot_23 = (|{_zz_PmpPlugin_logic_entries_2_napot_22,{_zz_PmpPlugin_logic_entries_2_napot_20,{_zz_PmpPlugin_logic_entries_2_napot_18,_zz_PmpPlugin_logic_entries_2_napot_17}}});
  assign PmpPlugin_logic_entries_2_napot = _zz_PmpPlugin_logic_entries_2_napot_24[20 : 1];
  always @(*) begin
    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_9 = (PmpPlugin_logic_entries_2_isNapot ? 10'h3ff : 10'h0);
    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_9[9] = (PmpPlugin_logic_entries_2_address[0] && PmpPlugin_logic_entries_2_isNapot);
  end

  always @(*) begin
    PmpPlugin_logic_entries_3_cfgNext_kind = PmpPlugin_logic_entries_3_cfg_kind;
    if(when_CsrAccessPlugin_l352_4) begin
      PmpPlugin_logic_entries_3_cfgNext_kind = CsrAccessPlugin_bus_write_bits[28 : 27];
    end
  end

  always @(*) begin
    PmpPlugin_logic_entries_3_cfgNext_read = PmpPlugin_logic_entries_3_cfg_read;
    if(when_CsrAccessPlugin_l352_4) begin
      PmpPlugin_logic_entries_3_cfgNext_read = CsrAccessPlugin_bus_write_bits[24];
    end
  end

  always @(*) begin
    PmpPlugin_logic_entries_3_cfgNext_write = PmpPlugin_logic_entries_3_cfg_write;
    if(when_CsrAccessPlugin_l352_4) begin
      PmpPlugin_logic_entries_3_cfgNext_write = CsrAccessPlugin_bus_write_bits[25];
    end
  end

  always @(*) begin
    PmpPlugin_logic_entries_3_cfgNext_execute = PmpPlugin_logic_entries_3_cfg_execute;
    if(when_CsrAccessPlugin_l352_4) begin
      PmpPlugin_logic_entries_3_cfgNext_execute = CsrAccessPlugin_bus_write_bits[26];
    end
  end

  always @(*) begin
    PmpPlugin_logic_entries_3_cfgNext_locked = PmpPlugin_logic_entries_3_cfg_locked;
    if(when_CsrAccessPlugin_l352_4) begin
      PmpPlugin_logic_entries_3_cfgNext_locked = CsrAccessPlugin_bus_write_bits[31];
    end
  end

  assign when_PmpPlugin_l127_3 = (! PmpPlugin_logic_entries_3_cfg_locked);
  assign when_PmpPlugin_l129_3 = (! PmpPlugin_logic_entries_3_cfgNext_read);
  assign _zz_PmpPlugin_logic_entries_3_napot = (~ PmpPlugin_logic_entries_3_address[19 : 0]);
  assign _zz_PmpPlugin_logic_entries_3_napot_1 = _zz_PmpPlugin_logic_entries_3_napot[0];
  assign _zz_PmpPlugin_logic_entries_3_napot_2 = _zz_PmpPlugin_logic_entries_3_napot[1];
  assign _zz_PmpPlugin_logic_entries_3_napot_3 = _zz_PmpPlugin_logic_entries_3_napot[2];
  assign _zz_PmpPlugin_logic_entries_3_napot_4 = _zz_PmpPlugin_logic_entries_3_napot[4];
  assign _zz_PmpPlugin_logic_entries_3_napot_5 = _zz_PmpPlugin_logic_entries_3_napot[5];
  assign _zz_PmpPlugin_logic_entries_3_napot_6 = _zz_PmpPlugin_logic_entries_3_napot[6];
  assign _zz_PmpPlugin_logic_entries_3_napot_7 = _zz_PmpPlugin_logic_entries_3_napot[8];
  assign _zz_PmpPlugin_logic_entries_3_napot_8 = _zz_PmpPlugin_logic_entries_3_napot[9];
  assign _zz_PmpPlugin_logic_entries_3_napot_9 = _zz_PmpPlugin_logic_entries_3_napot[10];
  assign _zz_PmpPlugin_logic_entries_3_napot_10 = _zz_PmpPlugin_logic_entries_3_napot[12];
  assign _zz_PmpPlugin_logic_entries_3_napot_11 = _zz_PmpPlugin_logic_entries_3_napot[13];
  assign _zz_PmpPlugin_logic_entries_3_napot_12 = _zz_PmpPlugin_logic_entries_3_napot[14];
  assign _zz_PmpPlugin_logic_entries_3_napot_13 = _zz_PmpPlugin_logic_entries_3_napot[16];
  assign _zz_PmpPlugin_logic_entries_3_napot_14 = _zz_PmpPlugin_logic_entries_3_napot[17];
  assign _zz_PmpPlugin_logic_entries_3_napot_15 = _zz_PmpPlugin_logic_entries_3_napot[18];
  always @(*) begin
    _zz_PmpPlugin_logic_entries_3_napot_16[0] = _zz_PmpPlugin_logic_entries_3_napot_1;
    _zz_PmpPlugin_logic_entries_3_napot_16[1] = (|{_zz_PmpPlugin_logic_entries_3_napot_2,_zz_PmpPlugin_logic_entries_3_napot_1});
    _zz_PmpPlugin_logic_entries_3_napot_16[2] = (|{_zz_PmpPlugin_logic_entries_3_napot_3,{_zz_PmpPlugin_logic_entries_3_napot_2,_zz_PmpPlugin_logic_entries_3_napot_1}});
    _zz_PmpPlugin_logic_entries_3_napot_16[3] = _zz_PmpPlugin_logic_entries_3_napot_17;
    _zz_PmpPlugin_logic_entries_3_napot_16[4] = (_zz_PmpPlugin_logic_entries_3_napot_4 || _zz_PmpPlugin_logic_entries_3_napot_17);
    _zz_PmpPlugin_logic_entries_3_napot_16[5] = ((|{_zz_PmpPlugin_logic_entries_3_napot_5,_zz_PmpPlugin_logic_entries_3_napot_4}) || _zz_PmpPlugin_logic_entries_3_napot_17);
    _zz_PmpPlugin_logic_entries_3_napot_16[6] = ((|{_zz_PmpPlugin_logic_entries_3_napot_6,{_zz_PmpPlugin_logic_entries_3_napot_5,_zz_PmpPlugin_logic_entries_3_napot_4}}) || _zz_PmpPlugin_logic_entries_3_napot_17);
    _zz_PmpPlugin_logic_entries_3_napot_16[7] = (_zz_PmpPlugin_logic_entries_3_napot_18 || _zz_PmpPlugin_logic_entries_3_napot_17);
    _zz_PmpPlugin_logic_entries_3_napot_16[8] = (_zz_PmpPlugin_logic_entries_3_napot_7 || _zz_PmpPlugin_logic_entries_3_napot_19);
    _zz_PmpPlugin_logic_entries_3_napot_16[9] = ((|{_zz_PmpPlugin_logic_entries_3_napot_8,_zz_PmpPlugin_logic_entries_3_napot_7}) || _zz_PmpPlugin_logic_entries_3_napot_19);
    _zz_PmpPlugin_logic_entries_3_napot_16[10] = ((|{_zz_PmpPlugin_logic_entries_3_napot_9,{_zz_PmpPlugin_logic_entries_3_napot_8,_zz_PmpPlugin_logic_entries_3_napot_7}}) || _zz_PmpPlugin_logic_entries_3_napot_19);
    _zz_PmpPlugin_logic_entries_3_napot_16[11] = (_zz_PmpPlugin_logic_entries_3_napot_20 || _zz_PmpPlugin_logic_entries_3_napot_19);
    _zz_PmpPlugin_logic_entries_3_napot_16[12] = (_zz_PmpPlugin_logic_entries_3_napot_10 || _zz_PmpPlugin_logic_entries_3_napot_21);
    _zz_PmpPlugin_logic_entries_3_napot_16[13] = ((|{_zz_PmpPlugin_logic_entries_3_napot_11,_zz_PmpPlugin_logic_entries_3_napot_10}) || _zz_PmpPlugin_logic_entries_3_napot_21);
    _zz_PmpPlugin_logic_entries_3_napot_16[14] = ((|{_zz_PmpPlugin_logic_entries_3_napot_12,{_zz_PmpPlugin_logic_entries_3_napot_11,_zz_PmpPlugin_logic_entries_3_napot_10}}) || _zz_PmpPlugin_logic_entries_3_napot_21);
    _zz_PmpPlugin_logic_entries_3_napot_16[15] = (_zz_PmpPlugin_logic_entries_3_napot_22 || _zz_PmpPlugin_logic_entries_3_napot_21);
    _zz_PmpPlugin_logic_entries_3_napot_16[16] = (_zz_PmpPlugin_logic_entries_3_napot_13 || _zz_PmpPlugin_logic_entries_3_napot_23);
    _zz_PmpPlugin_logic_entries_3_napot_16[17] = ((|{_zz_PmpPlugin_logic_entries_3_napot_14,_zz_PmpPlugin_logic_entries_3_napot_13}) || _zz_PmpPlugin_logic_entries_3_napot_23);
    _zz_PmpPlugin_logic_entries_3_napot_16[18] = ((|{_zz_PmpPlugin_logic_entries_3_napot_15,{_zz_PmpPlugin_logic_entries_3_napot_14,_zz_PmpPlugin_logic_entries_3_napot_13}}) || _zz_PmpPlugin_logic_entries_3_napot_23);
    _zz_PmpPlugin_logic_entries_3_napot_16[19] = ((|{_zz_PmpPlugin_logic_entries_3_napot[19],{_zz_PmpPlugin_logic_entries_3_napot_15,{_zz_PmpPlugin_logic_entries_3_napot_14,_zz_PmpPlugin_logic_entries_3_napot_13}}}) || _zz_PmpPlugin_logic_entries_3_napot_23);
  end

  assign _zz_PmpPlugin_logic_entries_3_napot_17 = (|{_zz_PmpPlugin_logic_entries_3_napot[3],{_zz_PmpPlugin_logic_entries_3_napot_3,{_zz_PmpPlugin_logic_entries_3_napot_2,_zz_PmpPlugin_logic_entries_3_napot_1}}});
  assign _zz_PmpPlugin_logic_entries_3_napot_18 = (|{_zz_PmpPlugin_logic_entries_3_napot[7],{_zz_PmpPlugin_logic_entries_3_napot_6,{_zz_PmpPlugin_logic_entries_3_napot_5,_zz_PmpPlugin_logic_entries_3_napot_4}}});
  assign _zz_PmpPlugin_logic_entries_3_napot_19 = (|{_zz_PmpPlugin_logic_entries_3_napot_18,_zz_PmpPlugin_logic_entries_3_napot_17});
  assign _zz_PmpPlugin_logic_entries_3_napot_20 = (|{_zz_PmpPlugin_logic_entries_3_napot[11],{_zz_PmpPlugin_logic_entries_3_napot_9,{_zz_PmpPlugin_logic_entries_3_napot_8,_zz_PmpPlugin_logic_entries_3_napot_7}}});
  assign _zz_PmpPlugin_logic_entries_3_napot_21 = (|{_zz_PmpPlugin_logic_entries_3_napot_20,{_zz_PmpPlugin_logic_entries_3_napot_18,_zz_PmpPlugin_logic_entries_3_napot_17}});
  assign _zz_PmpPlugin_logic_entries_3_napot_22 = (|{_zz_PmpPlugin_logic_entries_3_napot[15],{_zz_PmpPlugin_logic_entries_3_napot_12,{_zz_PmpPlugin_logic_entries_3_napot_11,_zz_PmpPlugin_logic_entries_3_napot_10}}});
  assign _zz_PmpPlugin_logic_entries_3_napot_23 = (|{_zz_PmpPlugin_logic_entries_3_napot_22,{_zz_PmpPlugin_logic_entries_3_napot_20,{_zz_PmpPlugin_logic_entries_3_napot_18,_zz_PmpPlugin_logic_entries_3_napot_17}}});
  assign PmpPlugin_logic_entries_3_napot = _zz_PmpPlugin_logic_entries_3_napot_24[20 : 1];
  always @(*) begin
    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_11 = (PmpPlugin_logic_entries_3_isNapot ? 10'h3ff : 10'h0);
    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_11[9] = (PmpPlugin_logic_entries_3_address[0] && PmpPlugin_logic_entries_3_isNapot);
  end

  assign PmpPlugin_logic_entries_0_isLocked = (PmpPlugin_logic_entries_0_cfg_locked || (PmpPlugin_logic_entries_1_cfg_locked && PmpPlugin_logic_entries_1_isTor));
  assign PmpPlugin_logic_entries_1_isLocked = (PmpPlugin_logic_entries_1_cfg_locked || (PmpPlugin_logic_entries_2_cfg_locked && PmpPlugin_logic_entries_2_isTor));
  assign PmpPlugin_logic_entries_2_isLocked = (PmpPlugin_logic_entries_2_cfg_locked || (PmpPlugin_logic_entries_3_cfg_locked && PmpPlugin_logic_entries_3_isTor));
  assign PmpPlugin_logic_entries_3_isLocked = (PmpPlugin_logic_entries_3_cfg_locked || 1'b0);
  always @(*) begin
    case(execute_ctrl2_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0)
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : begin
        early0_IntAluPlugin_logic_alu_bitwise = (execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0 & execute_ctrl2_down_early0_SrcPlugin_SRC2_lane0);
      end
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : begin
        early0_IntAluPlugin_logic_alu_bitwise = (execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0 | execute_ctrl2_down_early0_SrcPlugin_SRC2_lane0);
      end
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : begin
        early0_IntAluPlugin_logic_alu_bitwise = (execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0 ^ execute_ctrl2_down_early0_SrcPlugin_SRC2_lane0);
      end
      default : begin
        early0_IntAluPlugin_logic_alu_bitwise = 64'h0;
      end
    endcase
  end

  assign early0_IntAluPlugin_logic_alu_result = (_zz_early0_IntAluPlugin_logic_alu_result | _zz_early0_IntAluPlugin_logic_alu_result_2);
  assign execute_ctrl2_down_early0_IntAluPlugin_ALU_RESULT_lane0 = early0_IntAluPlugin_logic_alu_result;
  assign early0_IntAluPlugin_logic_wb_valid = execute_ctrl2_down_early0_IntAluPlugin_SEL_lane0;
  assign early0_IntAluPlugin_logic_wb_payload = execute_ctrl2_down_early0_IntAluPlugin_ALU_RESULT_lane0;
  always @(*) begin
    early0_BarrelShifterPlugin_logic_shift_amplitude = _zz_early0_BarrelShifterPlugin_logic_shift_amplitude;
    if(execute_ctrl2_down_BarrelShifterPlugin_IS_W_lane0) begin
      early0_BarrelShifterPlugin_logic_shift_amplitude[5] = 1'b0;
    end
  end

  always @(*) begin
    early0_BarrelShifterPlugin_logic_shift_reversed = (execute_ctrl2_down_BarrelShifterPlugin_LEFT_lane0 ? _zz_early0_BarrelShifterPlugin_logic_shift_reversed : execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0);
    if(execute_ctrl2_down_BarrelShifterPlugin_IS_W_RIGHT_lane0) begin
      early0_BarrelShifterPlugin_logic_shift_reversed[63 : 32] = ((execute_ctrl2_down_BarrelShifterPlugin_SIGNED_lane0 && execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[31]) ? 32'hffffffff : 32'h0);
    end
  end

  assign early0_BarrelShifterPlugin_logic_shift_shifted = _zz_early0_BarrelShifterPlugin_logic_shift_shifted[63:0];
  assign early0_BarrelShifterPlugin_logic_shift_patched = (execute_ctrl2_down_BarrelShifterPlugin_LEFT_lane0 ? _zz_early0_BarrelShifterPlugin_logic_shift_patched : early0_BarrelShifterPlugin_logic_shift_shifted);
  assign execute_ctrl2_down_early0_BarrelShifterPlugin_SHIFT_RESULT_lane0 = early0_BarrelShifterPlugin_logic_shift_patched;
  assign early0_BarrelShifterPlugin_logic_wb_valid = execute_ctrl2_down_early0_BarrelShifterPlugin_SEL_lane0;
  assign early0_BarrelShifterPlugin_logic_wb_payload = execute_ctrl2_down_early0_BarrelShifterPlugin_SHIFT_RESULT_lane0;
  always @(*) begin
    LsuPlugin_logic_events_waiting = 1'b0;
    if(LsuPlugin_logic_onCtrl_hartRegulation_valid) begin
      LsuPlugin_logic_events_waiting = 1'b1;
    end
  end

  always @(*) begin
    LsuL1_ackUnlock = 1'b0;
    if(LsuPlugin_logic_onCtrl_io_cmdSent) begin
      LsuL1_ackUnlock = 1'b1;
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_banksWrite_address = 9'bxxxxxxxxx;
    LsuL1Plugin_logic_banksWrite_address = {LsuL1Plugin_logic_refill_read_rspAddress[11 : 6],LsuL1Plugin_logic_refill_read_wordIndex};
    if(LsuL1Plugin_logic_lsu_ctrl_bankWriteReservation_win) begin
      LsuL1Plugin_logic_banksWrite_address = execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0[11 : 3];
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_banksWrite_writeData = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    LsuL1Plugin_logic_banksWrite_writeData = LsuL1Plugin_logic_bus_read_rsp_payload_data;
    if(LsuL1Plugin_logic_lsu_ctrl_bankWriteReservation_win) begin
      LsuL1Plugin_logic_banksWrite_writeData[63 : 0] = execute_ctrl4_down_LsuL1_WRITE_DATA_lane0;
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_banksWrite_writeMask = 8'bxxxxxxxx;
    LsuL1Plugin_logic_banksWrite_writeMask = 8'hff;
    if(LsuL1Plugin_logic_lsu_ctrl_bankWriteReservation_win) begin
      LsuL1Plugin_logic_banksWrite_writeMask = 8'h0;
      if(_zz_when[0]) begin
        LsuL1Plugin_logic_banksWrite_writeMask[7 : 0] = execute_ctrl4_down_LsuL1_MASK_lane0;
      end
    end
    if(LsuL1Plugin_logic_lsu_ctrl_preventSideEffects) begin
      if(LsuL1Plugin_logic_lsu_ctrl_bankWriteReservation_win) begin
        LsuL1Plugin_logic_banksWrite_writeMask = 8'h0;
      end
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_waysWrite_mask = 2'b00;
    if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
      if(when_LsuL1Plugin_l466) begin
        LsuL1Plugin_logic_waysWrite_mask[LsuL1Plugin_logic_refill_read_way] = 1'b1;
      end
    end
    if(LsuL1Plugin_logic_lsu_ctrl_doCbm) begin
      LsuL1Plugin_logic_waysWrite_mask = execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0;
    end
    if(LsuL1Plugin_logic_lsu_ctrl_doFlush) begin
      LsuL1Plugin_logic_waysWrite_mask = LsuL1Plugin_logic_lsu_ctrl_needFlushOh;
    end
    if(LsuL1Plugin_logic_lsu_ctrl_preventSideEffects) begin
      if(LsuL1Plugin_logic_lsu_ctrl_wayWriteReservation_win) begin
        LsuL1Plugin_logic_waysWrite_mask = 2'b00;
      end
    end
    if(when_LsuL1Plugin_l1233) begin
      LsuL1Plugin_logic_waysWrite_mask = 2'b11;
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_waysWrite_address = 6'bxxxxxx;
    if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
      if(when_LsuL1Plugin_l466) begin
        LsuL1Plugin_logic_waysWrite_address = LsuL1Plugin_logic_refill_read_rspAddress[11 : 6];
      end
    end
    if(LsuL1Plugin_logic_lsu_ctrl_doCbm) begin
      LsuL1Plugin_logic_waysWrite_address = execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0[11 : 6];
    end
    if(LsuL1Plugin_logic_lsu_ctrl_doFlush) begin
      LsuL1Plugin_logic_waysWrite_address = execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0[11 : 6];
    end
    if(when_LsuL1Plugin_l1233) begin
      LsuL1Plugin_logic_waysWrite_address = LsuL1Plugin_logic_initializer_counter[5:0];
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_waysWrite_tag_loaded = 1'bx;
    if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
      if(when_LsuL1Plugin_l466) begin
        LsuL1Plugin_logic_waysWrite_tag_loaded = 1'b1;
      end
    end
    if(LsuL1Plugin_logic_lsu_ctrl_doCbm) begin
      LsuL1Plugin_logic_waysWrite_tag_loaded = (! execute_ctrl4_down_LsuL1_INVALID_lane0);
    end
    if(LsuL1Plugin_logic_lsu_ctrl_doFlush) begin
      LsuL1Plugin_logic_waysWrite_tag_loaded = 1'b1;
    end
    if(when_LsuL1Plugin_l1233) begin
      LsuL1Plugin_logic_waysWrite_tag_loaded = 1'b0;
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_waysWrite_tag_address = 20'bxxxxxxxxxxxxxxxxxxxx;
    if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
      if(when_LsuL1Plugin_l466) begin
        LsuL1Plugin_logic_waysWrite_tag_address = LsuL1Plugin_logic_refill_read_rspAddress[31 : 12];
      end
    end
    if(LsuL1Plugin_logic_lsu_ctrl_doCbm) begin
      LsuL1Plugin_logic_waysWrite_tag_address = execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0[31 : 12];
    end
    if(LsuL1Plugin_logic_lsu_ctrl_doFlush) begin
      LsuL1Plugin_logic_waysWrite_tag_address = _zz_LsuL1Plugin_logic_waysWrite_tag_address;
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_waysWrite_tag_fault = 1'bx;
    if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
      if(when_LsuL1Plugin_l466) begin
        LsuL1Plugin_logic_waysWrite_tag_fault = LsuL1Plugin_logic_refill_read_faulty;
      end
    end
    if(LsuL1Plugin_logic_lsu_ctrl_doCbm) begin
      LsuL1Plugin_logic_waysWrite_tag_fault = _zz_LsuL1Plugin_logic_waysWrite_tag_fault[0];
    end
    if(LsuL1Plugin_logic_lsu_ctrl_doFlush) begin
      LsuL1Plugin_logic_waysWrite_tag_fault = _zz_LsuL1Plugin_logic_waysWrite_tag_fault_1;
    end
  end

  assign LsuL1Plugin_logic_waysWrite_valid = (|LsuL1Plugin_logic_waysWrite_mask);
  assign LsuL1Plugin_logic_banks_0_write_valid = LsuL1Plugin_logic_banksWrite_mask[0];
  assign LsuL1Plugin_logic_banks_0_write_payload_address = LsuL1Plugin_logic_banksWrite_address;
  assign LsuL1Plugin_logic_banks_0_write_payload_data = LsuL1Plugin_logic_banksWrite_writeData;
  assign LsuL1Plugin_logic_banks_0_write_payload_mask = LsuL1Plugin_logic_banksWrite_writeMask;
  assign LsuL1Plugin_logic_banks_0_read_rsp = LsuL1Plugin_logic_banks_0_mem_spinal_port1;
  assign LsuL1Plugin_logic_banks_1_write_valid = LsuL1Plugin_logic_banksWrite_mask[1];
  assign LsuL1Plugin_logic_banks_1_write_payload_address = LsuL1Plugin_logic_banksWrite_address;
  assign LsuL1Plugin_logic_banks_1_write_payload_data = LsuL1Plugin_logic_banksWrite_writeData;
  assign LsuL1Plugin_logic_banks_1_write_payload_mask = LsuL1Plugin_logic_banksWrite_writeMask;
  assign LsuL1Plugin_logic_banks_1_read_rsp = LsuL1Plugin_logic_banks_1_mem_spinal_port1;
  assign _zz_LsuL1Plugin_logic_ways_0_lsuRead_rsp_loaded = LsuL1Plugin_logic_ways_0_mem_spinal_port1;
  assign LsuL1Plugin_logic_ways_0_lsuRead_rsp_loaded = _zz_LsuL1Plugin_logic_ways_0_lsuRead_rsp_loaded[0];
  assign LsuL1Plugin_logic_ways_0_lsuRead_rsp_address = _zz_LsuL1Plugin_logic_ways_0_lsuRead_rsp_loaded[20 : 1];
  assign LsuL1Plugin_logic_ways_0_lsuRead_rsp_fault = _zz_LsuL1Plugin_logic_ways_0_lsuRead_rsp_loaded[21];
  assign _zz_LsuL1Plugin_logic_ways_1_lsuRead_rsp_loaded = LsuL1Plugin_logic_ways_1_mem_spinal_port1;
  assign LsuL1Plugin_logic_ways_1_lsuRead_rsp_loaded = _zz_LsuL1Plugin_logic_ways_1_lsuRead_rsp_loaded[0];
  assign LsuL1Plugin_logic_ways_1_lsuRead_rsp_address = _zz_LsuL1Plugin_logic_ways_1_lsuRead_rsp_loaded[20 : 1];
  assign LsuL1Plugin_logic_ways_1_lsuRead_rsp_fault = _zz_LsuL1Plugin_logic_ways_1_lsuRead_rsp_loaded[21];
  assign _zz_LsuL1Plugin_logic_shared_lsuRead_rsp_plru_0 = LsuL1Plugin_logic_shared_mem_spinal_port1;
  assign LsuL1Plugin_logic_shared_lsuRead_rsp_plru_0 = _zz_LsuL1Plugin_logic_shared_lsuRead_rsp_plru_0_1[0 : 0];
  assign LsuL1Plugin_logic_shared_lsuRead_rsp_dirty = _zz_LsuL1Plugin_logic_shared_lsuRead_rsp_plru_0[2 : 1];
  assign LsuL1Plugin_logic_slotsFreezeHazard = 1'b0;
  assign LsuL1Plugin_logic_slotsFreeze = (execute_freeze_valid && (! LsuL1Plugin_logic_slotsFreezeHazard));
  always @(*) begin
    LsuL1Plugin_logic_refill_slots_0_loadedSet = 1'b0;
    if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
      if(when_LsuL1Plugin_l466) begin
        LsuL1Plugin_logic_refill_slots_0_loadedSet = 1'b1;
      end
    end
  end

  assign LsuL1Plugin_logic_refill_slots_0_loadedDone = (LsuL1Plugin_logic_refill_slots_0_loadedCounter == 1'b1);
  assign LsuL1Plugin_logic_refill_slots_0_free = ((! LsuL1Plugin_logic_refill_slots_0_valid) && 1'b1);
  assign LsuL1Plugin_logic_refill_slots_0_fire = ((LsuL1Plugin_logic_refill_slots_0_valid && (! LsuL1Plugin_logic_slotsFreeze)) && LsuL1Plugin_logic_refill_slots_0_loadedDone);
  assign LsuL1Plugin_logic_refill_free = LsuL1Plugin_logic_refill_slots_0_free;
  assign LsuL1Plugin_logic_refill_full = (&(! LsuL1Plugin_logic_refill_slots_0_free));
  assign when_LsuL1Plugin_l382 = (LsuL1Plugin_logic_refill_push_valid && LsuL1Plugin_logic_refill_free[0]);
  assign when_LsuL1Plugin_l386 = LsuL1Plugin_logic_refill_free[0];
  assign LsuL1Plugin_logic_refill_read_arbiter_slotsWithId_0_0 = ((LsuL1Plugin_logic_refill_slots_0_valid && (! LsuL1Plugin_logic_refill_slots_0_cmdSent)) && (LsuL1Plugin_logic_refill_slots_0_victim == 1'b0));
  assign LsuL1Plugin_logic_refill_read_arbiter_hits = LsuL1Plugin_logic_refill_read_arbiter_slotsWithId_0_0;
  assign LsuL1Plugin_logic_refill_read_arbiter_hit = (|LsuL1Plugin_logic_refill_read_arbiter_hits);
  always @(*) begin
    LsuL1Plugin_logic_refill_read_arbiter_oh = (LsuL1Plugin_logic_refill_read_arbiter_hits & 1'b1);
    if(when_LsuL1Plugin_l303) begin
      LsuL1Plugin_logic_refill_read_arbiter_oh = LsuL1Plugin_logic_refill_read_arbiter_lock;
    end
  end

  assign when_LsuL1Plugin_l303 = (|LsuL1Plugin_logic_refill_read_arbiter_lock);
  assign LsuL1Plugin_logic_bus_read_cmd_fire = (LsuL1Plugin_logic_bus_read_cmd_valid && LsuL1Plugin_logic_bus_read_cmd_ready);
  assign LsuL1Plugin_logic_refill_read_cmdAddress = {LsuL1Plugin_logic_refill_slots_0_address[31 : 6],6'h0};
  assign LsuL1Plugin_logic_bus_read_cmd_valid = LsuL1Plugin_logic_refill_read_arbiter_hit;
  assign LsuL1Plugin_logic_bus_read_cmd_payload_address = LsuL1Plugin_logic_refill_read_cmdAddress;
  assign LsuL1Plugin_logic_refill_read_rspAddress = LsuL1Plugin_logic_refill_slots_0_address;
  assign LsuL1Plugin_logic_refill_read_way = LsuL1Plugin_logic_refill_slots_0_way;
  assign LsuL1Plugin_logic_refill_read_rspWithData = 1'b1;
  always @(*) begin
    LsuL1Plugin_logic_refill_read_writeReservation_take = 1'b0;
    if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
      LsuL1Plugin_logic_refill_read_writeReservation_take = 1'b1;
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_refill_read_bankWriteNotif[0] = ((LsuL1Plugin_logic_bus_read_rsp_valid && LsuL1Plugin_logic_refill_read_rspWithData) && (LsuL1Plugin_logic_refill_read_way == 1'b0));
    LsuL1Plugin_logic_refill_read_bankWriteNotif[1] = ((LsuL1Plugin_logic_bus_read_rsp_valid && LsuL1Plugin_logic_refill_read_rspWithData) && (LsuL1Plugin_logic_refill_read_way == 1'b1));
  end

  always @(*) begin
    LsuL1Plugin_logic_banksWrite_mask[0] = LsuL1Plugin_logic_refill_read_bankWriteNotif[0];
    LsuL1Plugin_logic_banksWrite_mask[1] = LsuL1Plugin_logic_refill_read_bankWriteNotif[1];
    if(LsuL1Plugin_logic_lsu_ctrl_bankWriteReservation_win) begin
      if(when_LsuL1Plugin_l940) begin
        LsuL1Plugin_logic_banksWrite_mask[0] = ((1'b0 == LsuL1Plugin_logic_lsu_ctrl_wayId) && LsuL1Plugin_logic_lsu_ctrl_doWrite);
      end
      if(when_LsuL1Plugin_l940_1) begin
        LsuL1Plugin_logic_banksWrite_mask[1] = ((1'b1 == LsuL1Plugin_logic_lsu_ctrl_wayId) && LsuL1Plugin_logic_lsu_ctrl_doWrite);
      end
    end
  end

  assign when_LsuL1Plugin_l453 = (LsuL1Plugin_logic_bus_read_rsp_valid && LsuL1Plugin_logic_bus_read_rsp_payload_error);
  always @(*) begin
    LsuL1Plugin_logic_refill_read_fire = 1'b0;
    if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
      if(when_LsuL1Plugin_l466) begin
        LsuL1Plugin_logic_refill_read_fire = 1'b1;
      end
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_refill_read_reservation_take = 1'b0;
    if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
      if(when_LsuL1Plugin_l466) begin
        LsuL1Plugin_logic_refill_read_reservation_take = 1'b1;
      end
    end
  end

  assign LsuL1Plugin_logic_refill_read_faulty = (LsuL1Plugin_logic_refill_read_hadError || LsuL1Plugin_logic_bus_read_rsp_payload_error);
  always @(*) begin
    LsuL1Plugin_logic_refillCompletions = 1'b0;
    if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
      if(when_LsuL1Plugin_l466) begin
        LsuL1Plugin_logic_refillCompletions[0] = 1'b1;
      end
    end
  end

  assign LsuL1Plugin_logic_bus_read_rsp_ready = 1'b1;
  assign when_LsuL1Plugin_l466 = ((LsuL1Plugin_logic_refill_read_wordIndex == 3'b111) || (! LsuL1Plugin_logic_refill_read_rspWithData));
  assign LsuL1_REFILL_BUSY = ((! LsuL1Plugin_logic_refill_slots_0_loaded) && (! LsuL1Plugin_logic_refill_slots_0_loadedSet));
  always @(*) begin
    LsuL1Plugin_logic_writeback_slots_0_fire = 1'b0;
    if(LsuL1Plugin_logic_bus_write_rsp_valid) begin
      LsuL1Plugin_logic_writeback_slots_0_fire = 1'b1;
    end
  end

  assign LsuL1Plugin_logic_writeback_slots_0_timer_done = (LsuL1Plugin_logic_writeback_slots_0_timer_counter == 1'b1);
  assign when_LsuL1Plugin_l533 = ((LsuL1Plugin_logic_writeback_slots_0_timer_done && (! LsuL1Plugin_logic_slotsFreeze)) && (LsuL1Plugin_logic_writeback_slots_0_fire || (! LsuL1Plugin_logic_writeback_slots_0_busy)));
  assign LsuL1Plugin_logic_writeback_slots_0_free = (! LsuL1Plugin_logic_writeback_slots_0_valid);
  assign LsuL1_WRITEBACK_BUSY = LsuL1Plugin_logic_writeback_slots_0_valid;
  assign LsuL1Plugin_logic_writebackBusy = (|LsuL1Plugin_logic_writeback_slots_0_valid);
  assign LsuL1Plugin_logic_writeback_free = LsuL1Plugin_logic_writeback_slots_0_free;
  assign LsuL1Plugin_logic_writeback_full = (&(! LsuL1Plugin_logic_writeback_slots_0_free));
  always @(*) begin
    LsuL1Plugin_logic_writeback_push_valid = 1'b0;
    if(LsuL1Plugin_logic_lsu_ctrl_doCbm) begin
      LsuL1Plugin_logic_writeback_push_valid = (execute_ctrl4_down_LsuL1_CLEAN_lane0 && LsuL1Plugin_logic_lsu_ctrl_wasDirty);
    end
    if(LsuL1Plugin_logic_lsu_ctrl_doFlush) begin
      LsuL1Plugin_logic_writeback_push_valid = 1'b1;
    end
    if(LsuL1Plugin_logic_lsu_ctrl_doRefill) begin
      LsuL1Plugin_logic_writeback_push_valid = LsuL1Plugin_logic_lsu_ctrl_refillWayNeedWriteback;
    end
    if(LsuL1Plugin_logic_lsu_ctrl_preventSideEffects) begin
      LsuL1Plugin_logic_writeback_push_valid = 1'b0;
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_writeback_push_payload_address = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(LsuL1Plugin_logic_lsu_ctrl_doCbm) begin
      LsuL1Plugin_logic_writeback_push_payload_address = ({6'd0,{execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0[31 : 12],execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0[11 : 6]}} <<< 3'd6);
    end
    if(LsuL1Plugin_logic_lsu_ctrl_doFlush) begin
      LsuL1Plugin_logic_writeback_push_payload_address = ({6'd0,{_zz_LsuL1Plugin_logic_waysWrite_tag_address,execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0[11 : 6]}} <<< 3'd6);
    end
    if(LsuL1Plugin_logic_lsu_ctrl_doRefill) begin
      LsuL1Plugin_logic_writeback_push_payload_address = ({6'd0,{_zz_LsuL1Plugin_logic_writeback_push_payload_address,execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0[11 : 6]}} <<< 3'd6);
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_writeback_push_payload_way = 1'bx;
    if(LsuL1Plugin_logic_lsu_ctrl_doCbm) begin
      LsuL1Plugin_logic_writeback_push_payload_way = LsuL1Plugin_logic_lsu_ctrl_wayId;
    end
    if(LsuL1Plugin_logic_lsu_ctrl_doFlush) begin
      LsuL1Plugin_logic_writeback_push_payload_way = LsuL1Plugin_logic_lsu_ctrl_needFlushSel;
    end
    if(LsuL1Plugin_logic_lsu_ctrl_doRefill) begin
      LsuL1Plugin_logic_writeback_push_payload_way = LsuL1Plugin_logic_lsu_ctrl_targetWay;
    end
  end

  assign when_LsuL1Plugin_l559 = (LsuL1Plugin_logic_writeback_free[0] && LsuL1Plugin_logic_writeback_push_valid);
  assign when_LsuL1Plugin_l564 = LsuL1Plugin_logic_writeback_free[0];
  assign LsuL1Plugin_logic_writeback_read_arbiter_slotsWithId_0_0 = (LsuL1Plugin_logic_writeback_slots_0_valid && (! LsuL1Plugin_logic_writeback_slots_0_readCmdDone));
  assign LsuL1Plugin_logic_writeback_read_arbiter_hits = LsuL1Plugin_logic_writeback_read_arbiter_slotsWithId_0_0;
  assign LsuL1Plugin_logic_writeback_read_arbiter_hit = (|LsuL1Plugin_logic_writeback_read_arbiter_hits);
  always @(*) begin
    LsuL1Plugin_logic_writeback_read_arbiter_oh = (LsuL1Plugin_logic_writeback_read_arbiter_hits & 1'b1);
    if(when_LsuL1Plugin_l303_1) begin
      LsuL1Plugin_logic_writeback_read_arbiter_oh = LsuL1Plugin_logic_writeback_read_arbiter_lock;
    end
  end

  assign when_LsuL1Plugin_l303_1 = (|LsuL1Plugin_logic_writeback_read_arbiter_lock);
  assign LsuL1Plugin_logic_writeback_read_address = LsuL1Plugin_logic_writeback_slots_0_address;
  assign LsuL1Plugin_logic_writeback_read_way = LsuL1Plugin_logic_writeback_slots_0_way;
  assign LsuL1Plugin_logic_writeback_read_slotRead_valid = LsuL1Plugin_logic_writeback_read_arbiter_hit;
  assign LsuL1Plugin_logic_writeback_read_slotRead_payload_wordIndex = LsuL1Plugin_logic_writeback_read_wordIndex;
  assign LsuL1Plugin_logic_writeback_read_slotRead_payload_way = LsuL1Plugin_logic_writeback_read_way;
  assign LsuL1Plugin_logic_writeback_read_slotRead_payload_last = (LsuL1Plugin_logic_writeback_read_wordIndex == 3'b111);
  assign when_LsuL1Plugin_l608 = (LsuL1Plugin_logic_writeback_read_slotRead_valid && LsuL1Plugin_logic_writeback_read_slotRead_payload_last);
  always @(*) begin
    LsuL1Plugin_logic_banks_0_read_cmd_valid = LsuL1Plugin_logic_banks_0_usedByWriteback;
    if(when_LsuL1Plugin_l721) begin
      LsuL1Plugin_logic_banks_0_read_cmd_valid = 1'b1;
    end
  end

  assign LsuL1Plugin_logic_banks_0_usedByWriteback = (LsuL1Plugin_logic_writeback_read_slotRead_valid && (LsuL1Plugin_logic_writeback_read_way == 1'b0));
  always @(*) begin
    LsuL1Plugin_logic_banks_0_read_cmd_payload = {LsuL1Plugin_logic_writeback_read_address[11 : 6],LsuL1Plugin_logic_writeback_read_wordIndex};
    if(when_LsuL1Plugin_l722) begin
      LsuL1Plugin_logic_banks_0_read_cmd_payload = LsuL1Plugin_logic_lsu_rb0_readAddress;
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_banks_1_read_cmd_valid = LsuL1Plugin_logic_banks_1_usedByWriteback;
    if(when_LsuL1Plugin_l721_1) begin
      LsuL1Plugin_logic_banks_1_read_cmd_valid = 1'b1;
    end
  end

  assign LsuL1Plugin_logic_banks_1_usedByWriteback = (LsuL1Plugin_logic_writeback_read_slotRead_valid && (LsuL1Plugin_logic_writeback_read_way == 1'b1));
  always @(*) begin
    LsuL1Plugin_logic_banks_1_read_cmd_payload = {LsuL1Plugin_logic_writeback_read_address[11 : 6],LsuL1Plugin_logic_writeback_read_wordIndex};
    if(when_LsuL1Plugin_l722_1) begin
      LsuL1Plugin_logic_banks_1_read_cmd_payload = LsuL1Plugin_logic_lsu_rb0_readAddress;
    end
  end

  assign LsuL1Plugin_logic_writeback_read_readedData = _zz_LsuL1Plugin_logic_writeback_read_readedData;
  assign LsuL1Plugin_logic_writeback_write_arbiter_slotsWithId_0_0 = ((LsuL1Plugin_logic_writeback_slots_0_valid && LsuL1Plugin_logic_writeback_slots_0_victimBufferReady) && (! LsuL1Plugin_logic_writeback_slots_0_writeCmdDone));
  assign LsuL1Plugin_logic_writeback_write_arbiter_hits = LsuL1Plugin_logic_writeback_write_arbiter_slotsWithId_0_0;
  assign LsuL1Plugin_logic_writeback_write_arbiter_hit = (|LsuL1Plugin_logic_writeback_write_arbiter_hits);
  always @(*) begin
    LsuL1Plugin_logic_writeback_write_arbiter_oh = (LsuL1Plugin_logic_writeback_write_arbiter_hits & 1'b1);
    if(when_LsuL1Plugin_l303_2) begin
      LsuL1Plugin_logic_writeback_write_arbiter_oh = LsuL1Plugin_logic_writeback_write_arbiter_lock;
    end
  end

  assign when_LsuL1Plugin_l303_2 = (|LsuL1Plugin_logic_writeback_write_arbiter_lock);
  assign LsuL1Plugin_logic_writeback_write_last = (LsuL1Plugin_logic_writeback_write_wordIndex == 3'b111);
  assign LsuL1Plugin_logic_writeback_write_bufferRead_valid = LsuL1Plugin_logic_writeback_write_arbiter_hit;
  assign LsuL1Plugin_logic_writeback_write_bufferRead_payload_last = LsuL1Plugin_logic_writeback_write_last;
  assign LsuL1Plugin_logic_writeback_write_bufferRead_payload_address = LsuL1Plugin_logic_writeback_slots_0_address;
  assign LsuL1Plugin_logic_writeback_write_bufferRead_fire = (LsuL1Plugin_logic_writeback_write_bufferRead_valid && LsuL1Plugin_logic_writeback_write_bufferRead_ready);
  assign when_LsuL1Plugin_l679 = (LsuL1Plugin_logic_writeback_write_bufferRead_fire && LsuL1Plugin_logic_writeback_write_last);
  always @(*) begin
    LsuL1Plugin_logic_writeback_write_bufferRead_ready = LsuL1Plugin_logic_writeback_write_cmd_ready;
    if(when_Stream_l477) begin
      LsuL1Plugin_logic_writeback_write_bufferRead_ready = 1'b1;
    end
  end

  assign when_Stream_l477 = (! LsuL1Plugin_logic_writeback_write_cmd_valid);
  assign LsuL1Plugin_logic_writeback_write_cmd_valid = LsuL1Plugin_logic_writeback_write_bufferRead_rValid;
  assign LsuL1Plugin_logic_writeback_write_cmd_payload_address = LsuL1Plugin_logic_writeback_write_bufferRead_rData_address;
  assign LsuL1Plugin_logic_writeback_write_cmd_payload_last = LsuL1Plugin_logic_writeback_write_bufferRead_rData_last;
  assign _zz_LsuL1Plugin_logic_writeback_write_word = LsuL1Plugin_logic_writeback_write_wordIndex;
  assign LsuL1Plugin_logic_writeback_write_word = LsuL1Plugin_logic_writeback_victimBuffer_spinal_port1;
  assign LsuL1Plugin_logic_bus_write_cmd_valid = LsuL1Plugin_logic_writeback_write_cmd_valid;
  assign LsuL1Plugin_logic_writeback_write_cmd_ready = LsuL1Plugin_logic_bus_write_cmd_ready;
  assign LsuL1Plugin_logic_bus_write_cmd_payload_fragment_address = LsuL1Plugin_logic_writeback_write_cmd_payload_address;
  assign LsuL1Plugin_logic_bus_write_cmd_payload_fragment_data = LsuL1Plugin_logic_writeback_write_word;
  assign LsuL1Plugin_logic_bus_write_cmd_payload_last = LsuL1Plugin_logic_writeback_write_cmd_payload_last;
  assign LsuL1Plugin_logic_lsu_rb0_readAddress = execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0[11 : 3];
  always @(*) begin
    execute_ctrl2_down_LsuL1Plugin_logic_BANK_BUSY_lane0[0] = LsuL1Plugin_logic_banks_0_usedByWriteback;
    execute_ctrl2_down_LsuL1Plugin_logic_BANK_BUSY_lane0[1] = LsuL1Plugin_logic_banks_1_usedByWriteback;
  end

  assign when_LsuL1Plugin_l721 = (! execute_freeze_valid);
  assign when_LsuL1Plugin_l722 = (! LsuL1Plugin_logic_banks_0_usedByWriteback);
  assign when_LsuL1Plugin_l721_1 = (! execute_freeze_valid);
  assign when_LsuL1Plugin_l722_1 = (! LsuL1Plugin_logic_banks_1_usedByWriteback);
  assign when_LsuL1Plugin_l738 = (! execute_freeze_valid);
  assign execute_ctrl3_down_LsuL1Plugin_logic_BANKS_WORDS_lane0_0 = LsuL1Plugin_logic_banks_0_read_rsp;
  always @(*) begin
    execute_ctrl3_down_LsuL1Plugin_logic_BANK_BUSY_REMAPPED_lane0[0] = (execute_ctrl3_down_LsuL1Plugin_logic_BANK_BUSY_lane0[1'b0] || LsuL1Plugin_logic_lsu_rb1_onBanks_0_busyReg);
    execute_ctrl3_down_LsuL1Plugin_logic_BANK_BUSY_REMAPPED_lane0[1] = (execute_ctrl3_down_LsuL1Plugin_logic_BANK_BUSY_lane0[1'b1] || LsuL1Plugin_logic_lsu_rb1_onBanks_1_busyReg);
  end

  assign when_LsuL1Plugin_l738_1 = (! execute_freeze_valid);
  assign execute_ctrl3_down_LsuL1Plugin_logic_BANKS_WORDS_lane0_1 = LsuL1Plugin_logic_banks_1_read_rsp;
  assign execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0 = execute_ctrl3_down_LsuL1Plugin_logic_BANKS_WORDS_lane0_0[63 : 0];
  assign execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1 = execute_ctrl3_down_LsuL1Plugin_logic_BANKS_WORDS_lane0_1[63 : 0];
  assign _zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0 = execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0[0];
  assign _zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0_1 = execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0[1];
  assign execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0 = ((_zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0 ? execute_ctrl4_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0 : 64'h0) | (_zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0_1 ? execute_ctrl4_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1 : 64'h0));
  always @(*) begin
    execute_ctrl3_down_LsuL1Plugin_logic_WRITE_TO_READ_HAZARDS_lane0[0] = ((execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_VALID_lane0 && (execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_ADDRESS_lane0[31 : 3] == execute_ctrl3_down_LsuL1_PHYSICAL_ADDRESS_lane0[31 : 3])) && 1'b1);
    execute_ctrl3_down_LsuL1Plugin_logic_WRITE_TO_READ_HAZARDS_lane0[1] = ((execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_VALID_lane0 && (execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_ADDRESS_lane0[31 : 3] == execute_ctrl3_down_LsuL1_PHYSICAL_ADDRESS_lane0[31 : 3])) && 1'b1);
  end

  assign execute_ctrl2_up_LsuL1Plugin_logic_FREEZE_HAZARD_lane0 = 1'b0;
  assign execute_ctrl3_LsuL1Plugin_logic_FREEZE_HAZARD_lane0_bypass = (execute_ctrl3_up_LsuL1Plugin_logic_FREEZE_HAZARD_lane0 || LsuL1Plugin_logic_slotsFreezeHazard);
  assign execute_ctrl4_LsuL1Plugin_logic_FREEZE_HAZARD_lane0_bypass = (execute_ctrl4_up_LsuL1Plugin_logic_FREEZE_HAZARD_lane0 || LsuL1Plugin_logic_slotsFreezeHazard);
  assign LsuL1Plugin_logic_shared_lsuRead_cmd_valid = (! execute_freeze_valid);
  assign LsuL1Plugin_logic_shared_lsuRead_cmd_payload = execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0[11 : 6];
  assign execute_ctrl2_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALID_lane0 = (LsuL1Plugin_logic_shared_write_valid && (LsuL1Plugin_logic_shared_write_payload_address == execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0[11 : 6]));
  assign execute_ctrl2_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_plru_0 = LsuL1Plugin_logic_shared_write_payload_data_plru_0;
  assign execute_ctrl2_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_dirty = LsuL1Plugin_logic_shared_write_payload_data_dirty;
  assign LsuL1Plugin_logic_ways_0_lsuRead_cmd_valid = (! execute_freeze_valid);
  assign LsuL1Plugin_logic_ways_0_lsuRead_cmd_payload = execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0[11 : 6];
  assign LsuL1Plugin_logic_ways_1_lsuRead_cmd_valid = (! execute_freeze_valid);
  assign LsuL1Plugin_logic_ways_1_lsuRead_cmd_payload = execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0[11 : 6];
  always @(*) begin
    execute_ctrl3_up_LsuL1Plugin_logic_SHARED_lane0_plru_0 = LsuL1Plugin_logic_shared_lsuRead_rsp_plru_0;
    if(execute_ctrl3_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALID_lane0) begin
      execute_ctrl3_up_LsuL1Plugin_logic_SHARED_lane0_plru_0 = execute_ctrl3_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_plru_0;
    end
  end

  always @(*) begin
    execute_ctrl3_up_LsuL1Plugin_logic_SHARED_lane0_dirty = LsuL1Plugin_logic_shared_lsuRead_rsp_dirty;
    if(execute_ctrl3_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALID_lane0) begin
      execute_ctrl3_up_LsuL1Plugin_logic_SHARED_lane0_dirty = execute_ctrl3_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_dirty;
    end
  end

  assign execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_loaded = LsuL1Plugin_logic_ways_0_lsuRead_rsp_loaded;
  assign execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_address = LsuL1Plugin_logic_ways_0_lsuRead_rsp_address;
  assign execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault = LsuL1Plugin_logic_ways_0_lsuRead_rsp_fault;
  assign execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_loaded = LsuL1Plugin_logic_ways_1_lsuRead_rsp_loaded;
  assign execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_address = LsuL1Plugin_logic_ways_1_lsuRead_rsp_address;
  assign execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault = LsuL1Plugin_logic_ways_1_lsuRead_rsp_fault;
  assign LsuL1Plugin_logic_lsu_sharedBypassers_0_hit = (LsuL1Plugin_logic_shared_write_valid && (LsuL1Plugin_logic_shared_write_payload_address == execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[11 : 6]));
  assign execute_ctrl3_LsuL1Plugin_logic_SHARED_lane0_bypass_plru_0 = (LsuL1Plugin_logic_lsu_sharedBypassers_0_hit ? LsuL1Plugin_logic_shared_write_payload_data_plru_0 : execute_ctrl3_up_LsuL1Plugin_logic_SHARED_lane0_plru_0);
  assign execute_ctrl3_LsuL1Plugin_logic_SHARED_lane0_bypass_dirty = (LsuL1Plugin_logic_lsu_sharedBypassers_0_hit ? LsuL1Plugin_logic_shared_write_payload_data_dirty : execute_ctrl3_up_LsuL1Plugin_logic_SHARED_lane0_dirty);
  always @(*) begin
    execute_ctrl3_down_LsuL1Plugin_logic_WAYS_HITS_lane0[0] = (execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_loaded && (execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_address == execute_ctrl3_down_LsuL1_PHYSICAL_ADDRESS_lane0[31 : 12]));
    execute_ctrl3_down_LsuL1Plugin_logic_WAYS_HITS_lane0[1] = (execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_loaded && (execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_address == execute_ctrl3_down_LsuL1_PHYSICAL_ADDRESS_lane0[31 : 12]));
  end

  assign execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HIT_lane0 = (|execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0);
  assign execute_ctrl4_down_LsuL1Plugin_logic_NEED_UNIQUE_lane0 = (execute_ctrl4_down_LsuL1_STORE_lane0 || execute_ctrl4_down_LsuL1_ATOMIC_lane0);
  assign LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_evict_logic_0_state = LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_context_state_0[0];
  assign LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_evict_sel_0 = (! LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_evict_logic_0_state);
  assign LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_evict_id = LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_evict_sel_0;
  assign LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_update_state_0[0] = LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_update_id[0];
  assign LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_context_state_0 = execute_ctrl4_down_LsuL1Plugin_logic_SHARED_lane0_plru_0;
  always @(*) begin
    LsuL1Plugin_logic_lsu_ctrl_wayWriteReservation_take = 1'b0;
    if(LsuL1Plugin_logic_lsu_ctrl_doCbm) begin
      LsuL1Plugin_logic_lsu_ctrl_wayWriteReservation_take = 1'b1;
    end
    if(LsuL1Plugin_logic_lsu_ctrl_doFlush) begin
      LsuL1Plugin_logic_lsu_ctrl_wayWriteReservation_take = 1'b1;
    end
  end

  assign LsuL1Plugin_logic_lsu_ctrl_bankWriteReservation_take = 1'b0;
  assign LsuL1Plugin_logic_lsu_ctrl_refillWayWithoutUpdate = LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_evict_id;
  assign LsuL1Plugin_logic_lsu_ctrl_refillWayNeedWriteback = _zz_LsuL1Plugin_logic_lsu_ctrl_refillWayNeedWriteback[LsuL1Plugin_logic_lsu_ctrl_refillWayWithoutUpdate];
  assign LsuL1Plugin_logic_lsu_ctrl_refillHazards = (LsuL1Plugin_logic_refill_slots_0_valid && (LsuL1Plugin_logic_refill_slots_0_address[11 : 6] == execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0[11 : 6]));
  assign LsuL1Plugin_logic_lsu_ctrl_writebackHazards = (LsuL1Plugin_logic_writeback_slots_0_valid && (LsuL1Plugin_logic_writeback_slots_0_address[11 : 6] == execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0[11 : 6]));
  assign LsuL1Plugin_logic_lsu_ctrl_refillHazard = (|LsuL1Plugin_logic_lsu_ctrl_refillHazards);
  assign LsuL1Plugin_logic_lsu_ctrl_writebackHazard = (|LsuL1Plugin_logic_lsu_ctrl_writebackHazards);
  assign LsuL1Plugin_logic_lsu_ctrl_wasDirty = (|(execute_ctrl4_down_LsuL1Plugin_logic_SHARED_lane0_dirty & execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0));
  assign LsuL1Plugin_logic_lsu_ctrl_loadedDirties = ({execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_loaded,execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_loaded} & execute_ctrl4_down_LsuL1Plugin_logic_SHARED_lane0_dirty);
  assign LsuL1Plugin_logic_lsu_ctrl_refillWayWasDirty = LsuL1Plugin_logic_lsu_ctrl_loadedDirties[LsuL1Plugin_logic_lsu_ctrl_refillWayWithoutUpdate];
  assign LsuL1Plugin_logic_lsu_ctrl_writeToReadHazard = 1'b0;
  assign LsuL1Plugin_logic_lsu_ctrl_bankNotRead = (|(execute_ctrl4_down_LsuL1Plugin_logic_BANK_BUSY_REMAPPED_lane0 & execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0));
  assign LsuL1Plugin_logic_lsu_ctrl_loadHazard = ((execute_ctrl4_down_LsuL1_LOAD_lane0 && (! execute_ctrl4_down_LsuL1_PREFETCH_lane0)) && (LsuL1Plugin_logic_lsu_ctrl_bankNotRead || LsuL1Plugin_logic_lsu_ctrl_writeToReadHazard));
  assign LsuL1Plugin_logic_lsu_ctrl_storeHazard = ((execute_ctrl4_down_LsuL1_STORE_lane0 && (! execute_ctrl4_down_LsuL1_PREFETCH_lane0)) && (! LsuL1Plugin_logic_lsu_ctrl_bankWriteReservation_win));
  assign LsuL1Plugin_logic_lsu_ctrl_preventSideEffects = (execute_ctrl4_down_LsuL1_ABORD_lane0 || execute_freeze_valid);
  assign LsuL1Plugin_logic_lsu_ctrl_flushHazard = (execute_ctrl4_down_LsuL1_FLUSH_lane0 && (! LsuL1Plugin_logic_lsu_ctrl_wayWriteReservation_win));
  assign LsuL1Plugin_logic_lsu_ctrl_coherencyHazard = 1'b0;
  assign execute_ctrl4_down_LsuL1Plugin_logic_HAZARD_FORCED_lane0 = 1'b0;
  assign execute_ctrl4_down_LsuL1_HAZARD_lane0 = ((((((LsuL1Plugin_logic_lsu_ctrl_hazardReg || LsuL1Plugin_logic_lsu_ctrl_loadHazard) || LsuL1Plugin_logic_lsu_ctrl_refillHazard) || LsuL1Plugin_logic_lsu_ctrl_storeHazard) || LsuL1Plugin_logic_lsu_ctrl_coherencyHazard) || execute_ctrl4_down_LsuL1Plugin_logic_HAZARD_FORCED_lane0) || execute_ctrl4_down_LsuL1Plugin_logic_FREEZE_HAZARD_lane0);
  assign execute_ctrl4_down_LsuL1_FLUSH_HAZARD_lane0 = (LsuL1Plugin_logic_lsu_ctrl_flushHazardReg || LsuL1Plugin_logic_lsu_ctrl_flushHazard);
  assign execute_ctrl4_down_LsuL1_MISS_lane0 = (! execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HIT_lane0);
  assign execute_ctrl4_down_LsuL1_FAULT_lane0 = ((execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HIT_lane0 && (|(execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0 & {execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault,execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault}))) && (! execute_ctrl4_down_LsuL1_FLUSH_lane0));
  assign execute_ctrl4_down_LsuL1_MISS_UNIQUE_lane0 = ((execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HIT_lane0 && execute_ctrl4_down_LsuL1Plugin_logic_NEED_UNIQUE_lane0) && 1'b0);
  assign execute_ctrl4_down_LsuL1_REFILL_HIT_lane0 = LsuL1Plugin_logic_lsu_ctrl_refillHazard;
  assign LsuL1Plugin_logic_events_loadAccess = ((((execute_ctrl4_up_LANE_SEL_lane0 && execute_ctrl4_up_isReady) && (! execute_lane0_ctrls_4_upIsCancel)) && execute_ctrl4_down_LsuL1_SEL_lane0) && execute_ctrl4_down_LsuL1_LOAD_lane0);
  assign LsuL1Plugin_logic_events_loadMiss = ((LsuL1Plugin_logic_events_loadAccess && (! execute_ctrl4_down_LsuL1_HAZARD_lane0)) && execute_ctrl4_down_LsuL1_MISS_lane0);
  assign LsuL1Plugin_logic_lsu_ctrl_canRefill = (((! (LsuL1Plugin_logic_lsu_ctrl_refillWayNeedWriteback && LsuL1Plugin_logic_writeback_full)) && (! LsuL1Plugin_logic_refill_full)) && (! LsuL1Plugin_logic_lsu_ctrl_writebackHazard));
  assign LsuL1Plugin_logic_lsu_ctrl_canFlush = (((LsuL1Plugin_logic_lsu_ctrl_wayWriteReservation_win && (! LsuL1Plugin_logic_writeback_full)) && (! (|LsuL1Plugin_logic_refill_slots_0_valid))) && (! LsuL1Plugin_logic_lsu_ctrl_writebackHazard));
  assign LsuL1Plugin_logic_lsu_ctrl_needFlushs = LsuL1Plugin_logic_lsu_ctrl_loadedDirties;
  assign _zz_LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_0 = LsuL1Plugin_logic_lsu_ctrl_needFlushs;
  assign LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_0 = _zz_LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_0[0];
  assign LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_1 = _zz_LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_0[1];
  always @(*) begin
    _zz_LsuL1Plugin_logic_lsu_ctrl_needFlushOh[0] = (LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_0 && (! 1'b0));
    _zz_LsuL1Plugin_logic_lsu_ctrl_needFlushOh[1] = (LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_1 && (! LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_0));
  end

  assign LsuL1Plugin_logic_lsu_ctrl_needFlushOh = _zz_LsuL1Plugin_logic_lsu_ctrl_needFlushOh;
  assign _zz_LsuL1Plugin_logic_lsu_ctrl_needFlushSel = LsuL1Plugin_logic_lsu_ctrl_needFlushOh[1];
  assign LsuL1Plugin_logic_lsu_ctrl_needFlushSel = _zz_LsuL1Plugin_logic_lsu_ctrl_needFlushSel;
  assign LsuL1Plugin_logic_lsu_ctrl_isAccess = ((! execute_ctrl4_down_LsuL1_FLUSH_lane0) && ((! execute_ctrl4_down_LsuL1_CLEAN_lane0) && (! execute_ctrl4_down_LsuL1_INVALID_lane0)));
  assign LsuL1Plugin_logic_lsu_ctrl_askRefill = ((LsuL1Plugin_logic_lsu_ctrl_isAccess && execute_ctrl4_down_LsuL1_MISS_lane0) && LsuL1Plugin_logic_lsu_ctrl_canRefill);
  assign LsuL1Plugin_logic_lsu_ctrl_askUpgrade = ((LsuL1Plugin_logic_lsu_ctrl_isAccess && execute_ctrl4_down_LsuL1_MISS_UNIQUE_lane0) && LsuL1Plugin_logic_lsu_ctrl_canRefill);
  assign LsuL1Plugin_logic_lsu_ctrl_askFlush = ((execute_ctrl4_down_LsuL1_FLUSH_lane0 && LsuL1Plugin_logic_lsu_ctrl_canFlush) && (|LsuL1Plugin_logic_lsu_ctrl_needFlushs));
  assign LsuL1Plugin_logic_lsu_ctrl_askCbm = (execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HIT_lane0 && (execute_ctrl4_down_LsuL1_INVALID_lane0 || (execute_ctrl4_down_LsuL1_CLEAN_lane0 && LsuL1Plugin_logic_lsu_ctrl_wasDirty)));
  assign LsuL1Plugin_logic_lsu_ctrl_doRefill = (execute_ctrl4_down_LsuL1_SEL_lane0 && LsuL1Plugin_logic_lsu_ctrl_askRefill);
  assign LsuL1Plugin_logic_lsu_ctrl_doUpgrade = (execute_ctrl4_down_LsuL1_SEL_lane0 && LsuL1Plugin_logic_lsu_ctrl_askUpgrade);
  assign LsuL1Plugin_logic_lsu_ctrl_doFlush = (execute_ctrl4_down_LsuL1_SEL_lane0 && LsuL1Plugin_logic_lsu_ctrl_askFlush);
  assign LsuL1Plugin_logic_lsu_ctrl_doWrite = ((((execute_ctrl4_down_LsuL1_SEL_lane0 && execute_ctrl4_down_LsuL1_STORE_lane0) && execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HIT_lane0) && _zz_LsuL1Plugin_logic_lsu_ctrl_doWrite[0]) && (! execute_ctrl4_down_LsuL1_SKIP_WRITE_lane0));
  assign LsuL1Plugin_logic_lsu_ctrl_doCbm = (((((execute_ctrl4_down_LsuL1_SEL_lane0 && LsuL1Plugin_logic_lsu_ctrl_askCbm) && LsuL1Plugin_logic_lsu_ctrl_wayWriteReservation_win) && (! LsuL1Plugin_logic_writeback_full)) && (! LsuL1Plugin_logic_lsu_ctrl_refillHazard)) && (! LsuL1Plugin_logic_lsu_ctrl_writebackHazard));
  assign LsuL1Plugin_logic_lsu_ctrl_wayId = _zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0_1;
  assign LsuL1Plugin_logic_lsu_ctrl_targetWay = (LsuL1Plugin_logic_lsu_ctrl_askUpgrade ? LsuL1Plugin_logic_lsu_ctrl_wayId : LsuL1Plugin_logic_lsu_ctrl_refillWayWithoutUpdate);
  always @(*) begin
    LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_update_id = LsuL1Plugin_logic_lsu_ctrl_wayId;
    if(LsuL1Plugin_logic_lsu_ctrl_doRefill) begin
      LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_update_id = LsuL1Plugin_logic_lsu_ctrl_targetWay;
    end
  end

  assign LsuL1Plugin_logic_lsu_ctrl_doRefillPush = (LsuL1Plugin_logic_lsu_ctrl_doRefill || LsuL1Plugin_logic_lsu_ctrl_doUpgrade);
  always @(*) begin
    LsuL1Plugin_logic_refill_push_valid = LsuL1Plugin_logic_lsu_ctrl_doRefillPush;
    if(LsuL1Plugin_logic_lsu_ctrl_preventSideEffects) begin
      LsuL1Plugin_logic_refill_push_valid = 1'b0;
    end
  end

  assign LsuL1Plugin_logic_refill_push_payload_address = execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0;
  assign LsuL1Plugin_logic_refill_push_payload_unique = execute_ctrl4_down_LsuL1Plugin_logic_NEED_UNIQUE_lane0;
  assign LsuL1Plugin_logic_refill_push_payload_data = LsuL1Plugin_logic_lsu_ctrl_askRefill;
  always @(*) begin
    LsuL1Plugin_logic_refill_push_payload_way = LsuL1Plugin_logic_lsu_ctrl_targetWay;
    if(LsuL1Plugin_logic_lsu_ctrl_askUpgrade) begin
      LsuL1Plugin_logic_refill_push_payload_way = LsuL1Plugin_logic_lsu_ctrl_wayId;
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_refill_push_payload_victim = ((LsuL1Plugin_logic_lsu_ctrl_refillWayNeedWriteback && LsuL1Plugin_logic_lsu_ctrl_refillWayWasDirty) ? LsuL1Plugin_logic_writeback_free : 1'b0);
    if(LsuL1Plugin_logic_lsu_ctrl_askUpgrade) begin
      LsuL1Plugin_logic_refill_push_payload_victim = 1'b0;
    end
  end

  assign execute_ctrl4_down_LsuL1_WAIT_REFILL_lane0 = (LsuL1Plugin_logic_lsu_ctrl_refillHazards | (((! execute_ctrl4_down_LsuL1_HAZARD_lane0) && (LsuL1Plugin_logic_lsu_ctrl_askRefill || LsuL1Plugin_logic_lsu_ctrl_askUpgrade)) ? (LsuL1Plugin_logic_refill_full ? 1'b1 : LsuL1Plugin_logic_refill_free) : 1'b0));
  assign execute_ctrl4_down_LsuL1_WAIT_WRITEBACK_lane0 = 1'b0;
  assign when_LsuL1Plugin_l926 = (execute_ctrl4_down_LsuL1_SEL_lane0 && (! execute_ctrl4_down_LsuL1_ABORD_lane0));
  assign _zz_22 = {LsuL1Plugin_logic_lsu_ctrl_askRefill,{LsuL1Plugin_logic_lsu_ctrl_doUpgrade,LsuL1Plugin_logic_lsu_ctrl_doFlush}};
  always @(*) begin
    LsuL1Plugin_logic_shared_write_valid = 1'b0;
    if(LsuL1Plugin_logic_lsu_ctrl_doCbm) begin
      LsuL1Plugin_logic_shared_write_valid = 1'b1;
    end
    if(LsuL1Plugin_logic_lsu_ctrl_doFlush) begin
      LsuL1Plugin_logic_shared_write_valid = 1'b1;
    end
    if(LsuL1Plugin_logic_lsu_ctrl_doRefill) begin
      LsuL1Plugin_logic_shared_write_valid = 1'b1;
    end
    if(when_LsuL1Plugin_l1028) begin
      LsuL1Plugin_logic_shared_write_valid = 1'b1;
    end
    if(LsuL1Plugin_logic_lsu_ctrl_preventSideEffects) begin
      LsuL1Plugin_logic_shared_write_valid = 1'b0;
    end
    if(when_LsuL1Plugin_l1233) begin
      LsuL1Plugin_logic_shared_write_valid = 1'b1;
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_shared_write_payload_address = execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0[11 : 6];
    if(when_LsuL1Plugin_l1233) begin
      LsuL1Plugin_logic_shared_write_payload_address = LsuL1Plugin_logic_initializer_counter[5:0];
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_shared_write_payload_data_plru_0 = LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_update_state_0;
    if(when_LsuL1Plugin_l1233) begin
      LsuL1Plugin_logic_shared_write_payload_data_plru_0 = _zz_LsuL1Plugin_logic_shared_write_payload_data_plru_0_1[0 : 0];
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_shared_write_payload_data_dirty = ((execute_ctrl4_down_LsuL1Plugin_logic_SHARED_lane0_dirty | (LsuL1Plugin_logic_lsu_ctrl_doWrite ? execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0 : 2'b00)) & (~ ((LsuL1Plugin_logic_lsu_ctrl_doRefill ? _zz_LsuL1Plugin_logic_shared_write_payload_data_dirty : 2'b00) | (LsuL1Plugin_logic_lsu_ctrl_doFlush ? LsuL1Plugin_logic_lsu_ctrl_needFlushOh : 2'b00))));
    if(LsuL1Plugin_logic_lsu_ctrl_doCbm) begin
      if(_zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0) begin
        LsuL1Plugin_logic_shared_write_payload_data_dirty[0] = 1'b0;
      end
      if(_zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0_1) begin
        LsuL1Plugin_logic_shared_write_payload_data_dirty[1] = 1'b0;
      end
    end
    if(when_LsuL1Plugin_l1233) begin
      LsuL1Plugin_logic_shared_write_payload_data_dirty = _zz_LsuL1Plugin_logic_shared_write_payload_data_plru_0[2 : 1];
    end
  end

  assign when_LsuL1Plugin_l940 = execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0[0];
  assign when_LsuL1Plugin_l940_1 = execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0[1];
  assign execute_ctrl4_down_LsuL1_CBM_REDO_lane0 = LsuL1Plugin_logic_lsu_ctrl_askCbm;
  assign execute_ctrl4_down_LsuL1_FLUSH_HIT_lane0 = (|LsuL1Plugin_logic_lsu_ctrl_needFlushs);
  assign _zz_LsuL1Plugin_logic_waysWrite_tag_address = _zz__zz_LsuL1Plugin_logic_waysWrite_tag_address;
  assign execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_VALID_lane0 = LsuL1Plugin_logic_lsu_ctrl_doWrite;
  assign execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_ADDRESS_lane0 = execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0;
  assign execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0 = execute_ctrl4_down_LsuL1_WRITE_DATA_lane0;
  assign execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0 = execute_ctrl4_down_LsuL1_MASK_lane0;
  assign when_LsuL1Plugin_l1028 = ((execute_ctrl4_down_LsuL1_SEL_lane0 && (! execute_ctrl4_down_LsuL1_HAZARD_lane0)) && (! execute_ctrl4_down_LsuL1_MISS_lane0));
  always @(*) begin
    execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0 = execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0;
    if(when_LsuL1Plugin_l1035) begin
      if(when_LsuL1Plugin_l1039) begin
        execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[7 : 0] = execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[7 : 0];
      end
      if(when_LsuL1Plugin_l1039_1) begin
        execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[15 : 8] = execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[15 : 8];
      end
      if(when_LsuL1Plugin_l1039_2) begin
        execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[23 : 16] = execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[23 : 16];
      end
      if(when_LsuL1Plugin_l1039_3) begin
        execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[31 : 24] = execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[31 : 24];
      end
      if(when_LsuL1Plugin_l1039_4) begin
        execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[39 : 32] = execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[39 : 32];
      end
      if(when_LsuL1Plugin_l1039_5) begin
        execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[47 : 40] = execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[47 : 40];
      end
      if(when_LsuL1Plugin_l1039_6) begin
        execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[55 : 48] = execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[55 : 48];
      end
      if(when_LsuL1Plugin_l1039_7) begin
        execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[63 : 56] = execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[63 : 56];
      end
    end
    if(when_LsuL1Plugin_l1035_1) begin
      if(when_LsuL1Plugin_l1039_8) begin
        execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[7 : 0] = execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[7 : 0];
      end
      if(when_LsuL1Plugin_l1039_9) begin
        execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[15 : 8] = execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[15 : 8];
      end
      if(when_LsuL1Plugin_l1039_10) begin
        execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[23 : 16] = execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[23 : 16];
      end
      if(when_LsuL1Plugin_l1039_11) begin
        execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[31 : 24] = execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[31 : 24];
      end
      if(when_LsuL1Plugin_l1039_12) begin
        execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[39 : 32] = execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[39 : 32];
      end
      if(when_LsuL1Plugin_l1039_13) begin
        execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[47 : 40] = execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[47 : 40];
      end
      if(when_LsuL1Plugin_l1039_14) begin
        execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[55 : 48] = execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[55 : 48];
      end
      if(when_LsuL1Plugin_l1039_15) begin
        execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[63 : 56] = execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[63 : 56];
      end
    end
  end

  assign when_LsuL1Plugin_l1035 = execute_ctrl4_down_LsuL1Plugin_logic_WRITE_TO_READ_HAZARDS_lane0[1];
  assign when_LsuL1Plugin_l1039 = execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[0];
  assign when_LsuL1Plugin_l1039_1 = execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[1];
  assign when_LsuL1Plugin_l1039_2 = execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[2];
  assign when_LsuL1Plugin_l1039_3 = execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[3];
  assign when_LsuL1Plugin_l1039_4 = execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[4];
  assign when_LsuL1Plugin_l1039_5 = execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[5];
  assign when_LsuL1Plugin_l1039_6 = execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[6];
  assign when_LsuL1Plugin_l1039_7 = execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[7];
  assign when_LsuL1Plugin_l1035_1 = execute_ctrl4_down_LsuL1Plugin_logic_WRITE_TO_READ_HAZARDS_lane0[0];
  assign when_LsuL1Plugin_l1039_8 = execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[0];
  assign when_LsuL1Plugin_l1039_9 = execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[1];
  assign when_LsuL1Plugin_l1039_10 = execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[2];
  assign when_LsuL1Plugin_l1039_11 = execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[3];
  assign when_LsuL1Plugin_l1039_12 = execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[4];
  assign when_LsuL1Plugin_l1039_13 = execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[5];
  assign when_LsuL1Plugin_l1039_14 = execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[6];
  assign when_LsuL1Plugin_l1039_15 = execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[7];
  assign execute_ctrl4_down_LsuL1_READ_DATA_lane0 = execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0;
  assign LsuL1Plugin_logic_initializer_done = LsuL1Plugin_logic_initializer_counter[6];
  assign when_LsuL1Plugin_l1233 = (! LsuL1Plugin_logic_initializer_done);
  assign _zz_LsuL1Plugin_logic_shared_write_payload_data_plru_0 = 3'b000;
  assign LsuL1Plugin_logic_refill_read_reservation_win = (! 1'b0);
  assign LsuL1Plugin_logic_lsu_ctrl_wayWriteReservation_win = (! (|LsuL1Plugin_logic_refill_read_reservation_take));
  assign LsuL1Plugin_logic_refill_read_writeReservation_win = (! 1'b0);
  assign LsuL1Plugin_logic_lsu_ctrl_bankWriteReservation_win = (! (|LsuL1Plugin_logic_refill_read_writeReservation_take));
  assign execute_ctrl2_down_MUL_SRC1_lane0 = _zz_execute_ctrl2_down_MUL_SRC1_lane0;
  assign execute_ctrl2_down_MUL_SRC2_lane0 = _zz_execute_ctrl2_down_MUL_SRC2_lane0;
  assign execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_0_lane0 = (execute_ctrl2_down_MUL_SRC1_lane0[16 : 0] * execute_ctrl2_down_MUL_SRC2_lane0[16 : 0]);
  assign execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_1_lane0 = (execute_ctrl2_down_MUL_SRC1_lane0[16 : 0] * execute_ctrl2_down_MUL_SRC2_lane0[33 : 17]);
  assign execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_2_lane0 = (execute_ctrl2_down_MUL_SRC1_lane0[33 : 17] * execute_ctrl2_down_MUL_SRC2_lane0[16 : 0]);
  assign execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_3_lane0 = (execute_ctrl2_down_MUL_SRC1_lane0[16 : 0] * execute_ctrl2_down_MUL_SRC2_lane0[50 : 34]);
  assign execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_4_lane0 = (execute_ctrl2_down_MUL_SRC1_lane0[33 : 17] * execute_ctrl2_down_MUL_SRC2_lane0[33 : 17]);
  assign execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_5_lane0 = (execute_ctrl2_down_MUL_SRC1_lane0[50 : 34] * execute_ctrl2_down_MUL_SRC2_lane0[16 : 0]);
  assign execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_6_lane0 = _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_6_lane0;
  assign execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_7_lane0 = _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_7_lane0;
  assign execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_8_lane0 = (execute_ctrl2_down_MUL_SRC1_lane0[33 : 17] * execute_ctrl2_down_MUL_SRC2_lane0[50 : 34]);
  assign execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_9_lane0 = (execute_ctrl2_down_MUL_SRC1_lane0[50 : 34] * execute_ctrl2_down_MUL_SRC2_lane0[33 : 17]);
  assign execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_10_lane0 = _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_10_lane0;
  assign execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_11_lane0 = _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_11_lane0;
  assign execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_12_lane0 = (execute_ctrl2_down_MUL_SRC1_lane0[50 : 34] * execute_ctrl2_down_MUL_SRC2_lane0[50 : 34]);
  assign execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_13_lane0 = _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_13_lane0;
  assign execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_14_lane0 = _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_14_lane0;
  assign execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_15_lane0 = _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_15_lane0;
  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0 = 61'h0;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0[33 : 0] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_0_lane0[33 : 0];
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0[60 : 34] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_3_lane0[26 : 0];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_1 = 61'h0;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_1[50 : 17] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_1_lane0[33 : 0];
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_1[60 : 51] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_6_lane0[9 : 0];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_2 = 61'h0;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_2[50 : 17] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_2_lane0[33 : 0];
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_2[60 : 51] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_7_lane0[9 : 0];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_3 = 61'h0;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_3[60 : 34] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_4_lane0[26 : 0];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_4 = 61'h0;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_4[60 : 34] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_5_lane0[26 : 0];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_5 = 61'h0;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_5[60 : 51] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_8_lane0[9 : 0];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_6 = 61'h0;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_6[60 : 51] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_9_lane0[9 : 0];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0 = 44'h0;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0[6 : 0] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_3_lane0[33 : 27];
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0[43 : 7] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_10_lane0[36 : 0];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_1 = 44'h0;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_1[43 : 0] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_6_lane0[53 : 10];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_2 = 44'h0;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_2[43 : 0] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_7_lane0[53 : 10];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_3 = 44'h0;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_3[6 : 0] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_4_lane0[33 : 27];
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_3[43 : 7] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_11_lane0[36 : 0];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_4 = 44'h0;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_4[6 : 0] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_5_lane0[33 : 27];
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_4[40 : 7] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_12_lane0[33 : 0];
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_4[43 : 41] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_15_lane0[2 : 0];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_5 = 44'h0;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_5[23 : 0] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_8_lane0[33 : 10];
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_5[43 : 24] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_13_lane0[19 : 0];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_6 = 44'h0;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_6[23 : 0] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_9_lane0[33 : 10];
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_6[43 : 24] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_14_lane0[19 : 0];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0 = 23'h0;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0[22 : 0] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_10_lane0[59 : 37];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_1 = 23'h0;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_1[22 : 0] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_6_lane0[76 : 54];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_2 = 23'h0;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_2[22 : 0] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_7_lane0[76 : 54];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_3 = 23'h0;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_3[22 : 0] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_11_lane0[59 : 37];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_4 = 23'h0;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_4[22 : 0] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_15_lane0[25 : 3];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_5 = 23'h0;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_5[22 : 0] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_13_lane0[42 : 20];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_6 = 23'h0;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_6[22 : 0] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_14_lane0[42 : 20];
  end

  assign execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0 = (_zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_7 + _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_14);
  assign execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0 = (_zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_7 + _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_14);
  assign execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0 = (_zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_7 + _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_14);
  always @(*) begin
    _zz_execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0 = 131'h0;
    _zz_execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0[63 : 0] = execute_ctrl4_down_early0_MulPlugin_logic_steps_0_adders_0_lane0[63 : 0];
    _zz_execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0[130 : 105] = execute_ctrl4_down_early0_MulPlugin_logic_steps_0_adders_2_lane0[25 : 0];
  end

  always @(*) begin
    _zz_execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0_1 = 131'h0;
    _zz_execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0_1[107 : 61] = execute_ctrl4_down_early0_MulPlugin_logic_steps_0_adders_1_lane0[46 : 0];
  end

  assign execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0 = (_zz_execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0 + _zz_execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0_1);
  assign early0_MulPlugin_logic_formatBus_valid = execute_ctrl4_down_early0_MulPlugin_SEL_lane0;
  assign early0_MulPlugin_logic_formatBus_payload = (execute_ctrl4_down_MulPlugin_HIGH_lane0 ? early0_MulPlugin_logic_writeback_buffer_data : execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0[63 : 0]);
  always @(*) begin
    execute_ctrl2_down_RsUnsignedPlugin_RS1_FORMATED_lane0 = execute_ctrl2_up_integer_RS1_lane0;
    if(execute_ctrl2_down_RsUnsignedPlugin_IS_W_lane0) begin
      execute_ctrl2_down_RsUnsignedPlugin_RS1_FORMATED_lane0[63 : 32] = ((execute_ctrl2_down_RsUnsignedPlugin_RS1_SIGNED_lane0 && execute_ctrl2_up_integer_RS1_lane0[31]) ? 32'hffffffff : 32'h0);
    end
  end

  always @(*) begin
    execute_ctrl2_down_RsUnsignedPlugin_RS2_FORMATED_lane0 = execute_ctrl2_up_integer_RS2_lane0;
    if(execute_ctrl2_down_RsUnsignedPlugin_IS_W_lane0) begin
      execute_ctrl2_down_RsUnsignedPlugin_RS2_FORMATED_lane0[63 : 32] = ((execute_ctrl2_down_RsUnsignedPlugin_RS2_SIGNED_lane0 && execute_ctrl2_up_integer_RS2_lane0[31]) ? 32'hffffffff : 32'h0);
    end
  end

  assign execute_ctrl2_down_RsUnsignedPlugin_RS1_REVERT_lane0 = (execute_ctrl2_down_RsUnsignedPlugin_RS1_SIGNED_lane0 && execute_ctrl2_down_RsUnsignedPlugin_RS1_FORMATED_lane0[63]);
  assign execute_ctrl2_down_RsUnsignedPlugin_RS2_REVERT_lane0 = (execute_ctrl2_down_RsUnsignedPlugin_RS2_SIGNED_lane0 && execute_ctrl2_down_RsUnsignedPlugin_RS2_FORMATED_lane0[63]);
  assign execute_ctrl2_down_RsUnsignedPlugin_RS1_UNSIGNED_lane0 = ((execute_ctrl2_down_RsUnsignedPlugin_RS1_REVERT_lane0 ? (~ execute_ctrl2_down_RsUnsignedPlugin_RS1_FORMATED_lane0) : execute_ctrl2_down_RsUnsignedPlugin_RS1_FORMATED_lane0) + _zz_execute_ctrl2_down_RsUnsignedPlugin_RS1_UNSIGNED_lane0);
  assign execute_ctrl2_down_RsUnsignedPlugin_RS2_UNSIGNED_lane0 = ((execute_ctrl2_down_RsUnsignedPlugin_RS2_REVERT_lane0 ? (~ execute_ctrl2_down_RsUnsignedPlugin_RS2_FORMATED_lane0) : execute_ctrl2_down_RsUnsignedPlugin_RS2_FORMATED_lane0) + _zz_execute_ctrl2_down_RsUnsignedPlugin_RS2_UNSIGNED_lane0);
  assign io_cmd_fire = (early0_DivPlugin_logic_processing_div_io_cmd_valid && early0_DivPlugin_logic_processing_div_io_cmd_ready);
  assign early0_DivPlugin_logic_processing_request = (execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_down_early0_DivPlugin_SEL_lane0);
  assign early0_DivPlugin_logic_processing_a = execute_ctrl2_down_RsUnsignedPlugin_RS1_UNSIGNED_lane0;
  assign early0_DivPlugin_logic_processing_b = execute_ctrl2_down_RsUnsignedPlugin_RS2_UNSIGNED_lane0;
  always @(*) begin
    early0_DivPlugin_logic_processing_div_io_cmd_valid = (early0_DivPlugin_logic_processing_request && (! early0_DivPlugin_logic_processing_cmdSent));
    if(when_DivPlugin_l121) begin
      early0_DivPlugin_logic_processing_div_io_cmd_valid = 1'b0;
    end
  end

  assign when_DivPlugin_l121 = (! early0_DivPlugin_logic_processing_relaxer_hadRequest);
  assign early0_DivPlugin_logic_processing_freeze = ((early0_DivPlugin_logic_processing_request && (! early0_DivPlugin_logic_processing_div_io_rsp_valid)) && (! early0_DivPlugin_logic_processing_unscheduleRequest));
  assign early0_DivPlugin_logic_processing_selected = (execute_ctrl2_down_DivPlugin_REM_lane0 ? early0_DivPlugin_logic_processing_div_io_rsp_payload_remain : early0_DivPlugin_logic_processing_div_io_rsp_payload_result);
  assign _zz_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0 = early0_DivPlugin_logic_processing_selected;
  assign execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0 = _zz_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0_1;
  assign early0_DivPlugin_logic_formatBus_valid = execute_ctrl3_down_early0_DivPlugin_SEL_lane0;
  assign early0_DivPlugin_logic_formatBus_payload = execute_ctrl3_down_DivPlugin_DIV_RESULT_lane0;
  assign WhiteboxerPlugin_logic_fetch_fire = fetch_logic_ctrls_0_down_isFiring;
  assign PrivilegedPlugin_api_harts_0_allowInterrupts = 1'b1;
  assign PrivilegedPlugin_api_harts_0_allowException = 1'b1;
  assign PrivilegedPlugin_api_harts_0_allowEbreakException = 1'b1;
  assign PrivilegedPlugin_api_harts_0_fpuEnable = 1'b0;
  assign LsuL1Axi4Plugin_logic_axi_ar_valid = LsuL1Plugin_logic_bus_read_cmd_valid;
  assign LsuL1Axi4Plugin_logic_axi_ar_payload_addr = LsuL1Plugin_logic_bus_read_cmd_payload_address;
  assign LsuL1Axi4Plugin_logic_axi_ar_payload_cache = 4'b1111;
  assign LsuL1Axi4Plugin_logic_axi_ar_payload_prot = 3'b010;
  assign LsuL1Axi4Plugin_logic_axi_ar_payload_len = 8'h07;
  assign LsuL1Axi4Plugin_logic_axi_ar_payload_size = 3'b011;
  assign LsuL1Axi4Plugin_logic_axi_ar_payload_burst = 2'b01;
  assign LsuL1Plugin_logic_bus_read_cmd_ready = LsuL1Axi4Plugin_logic_axi_ar_ready;
  assign LsuL1Plugin_logic_bus_read_rsp_valid = LsuL1Axi4Plugin_logic_axi_r_valid;
  assign LsuL1Plugin_logic_bus_read_rsp_payload_data = LsuL1Axi4Plugin_logic_axi_r_payload_data;
  assign LsuL1Plugin_logic_bus_read_rsp_payload_error = (! (LsuL1Axi4Plugin_logic_axi_r_payload_resp == 2'b00));
  assign LsuL1Axi4Plugin_logic_axi_r_ready = 1'b1;
  always @(*) begin
    LsuL1Plugin_logic_bus_write_cmd_ready = 1'b1;
    if(when_Stream_l1253) begin
      LsuL1Plugin_logic_bus_write_cmd_ready = 1'b0;
    end
    if(when_Stream_l1253_1) begin
      LsuL1Plugin_logic_bus_write_cmd_ready = 1'b0;
    end
  end

  assign when_Stream_l1253 = ((! LsuL1Plugin_logic_bus_toAxi4_awRaw_ready) && LsuL1Plugin_logic_bus_write_cmd_fork2_logic_linkEnable_0);
  assign when_Stream_l1253_1 = ((! LsuL1Plugin_logic_bus_toAxi4_wRaw_ready) && LsuL1Plugin_logic_bus_write_cmd_fork2_logic_linkEnable_1);
  assign LsuL1Plugin_logic_bus_toAxi4_awRaw_valid = (LsuL1Plugin_logic_bus_write_cmd_valid && LsuL1Plugin_logic_bus_write_cmd_fork2_logic_linkEnable_0);
  assign LsuL1Plugin_logic_bus_toAxi4_awRaw_payload_last = LsuL1Plugin_logic_bus_write_cmd_payload_last;
  assign LsuL1Plugin_logic_bus_toAxi4_awRaw_payload_fragment_address = LsuL1Plugin_logic_bus_write_cmd_payload_fragment_address;
  assign LsuL1Plugin_logic_bus_toAxi4_awRaw_payload_fragment_data = LsuL1Plugin_logic_bus_write_cmd_payload_fragment_data;
  assign LsuL1Plugin_logic_bus_toAxi4_awRaw_fire = (LsuL1Plugin_logic_bus_toAxi4_awRaw_valid && LsuL1Plugin_logic_bus_toAxi4_awRaw_ready);
  assign LsuL1Plugin_logic_bus_toAxi4_wRaw_valid = (LsuL1Plugin_logic_bus_write_cmd_valid && LsuL1Plugin_logic_bus_write_cmd_fork2_logic_linkEnable_1);
  assign LsuL1Plugin_logic_bus_toAxi4_wRaw_payload_last = LsuL1Plugin_logic_bus_write_cmd_payload_last;
  assign LsuL1Plugin_logic_bus_toAxi4_wRaw_payload_fragment_address = LsuL1Plugin_logic_bus_write_cmd_payload_fragment_address;
  assign LsuL1Plugin_logic_bus_toAxi4_wRaw_payload_fragment_data = LsuL1Plugin_logic_bus_write_cmd_payload_fragment_data;
  assign LsuL1Plugin_logic_bus_toAxi4_wRaw_fire = (LsuL1Plugin_logic_bus_toAxi4_wRaw_valid && LsuL1Plugin_logic_bus_toAxi4_wRaw_ready);
  assign when_Stream_l581 = (! LsuL1Plugin_logic_bus_toAxi4_awRaw_payload_first);
  always @(*) begin
    LsuL1Plugin_logic_bus_toAxi4_awFiltred_valid = LsuL1Plugin_logic_bus_toAxi4_awRaw_valid;
    if(when_Stream_l581) begin
      LsuL1Plugin_logic_bus_toAxi4_awFiltred_valid = 1'b0;
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_bus_toAxi4_awRaw_ready = LsuL1Plugin_logic_bus_toAxi4_awFiltred_ready;
    if(when_Stream_l581) begin
      LsuL1Plugin_logic_bus_toAxi4_awRaw_ready = 1'b1;
    end
  end

  assign LsuL1Plugin_logic_bus_toAxi4_awFiltred_payload_last = LsuL1Plugin_logic_bus_toAxi4_awRaw_payload_last;
  assign LsuL1Plugin_logic_bus_toAxi4_awFiltred_payload_fragment_address = LsuL1Plugin_logic_bus_toAxi4_awRaw_payload_fragment_address;
  assign LsuL1Plugin_logic_bus_toAxi4_awFiltred_payload_fragment_data = LsuL1Plugin_logic_bus_toAxi4_awRaw_payload_fragment_data;
  always @(*) begin
    LsuL1Plugin_logic_bus_toAxi4_awFiltred_ready = LsuL1Plugin_logic_bus_toAxi4_aw_ready;
    if(when_Stream_l477_1) begin
      LsuL1Plugin_logic_bus_toAxi4_awFiltred_ready = 1'b1;
    end
  end

  assign when_Stream_l477_1 = (! LsuL1Plugin_logic_bus_toAxi4_aw_valid);
  assign LsuL1Plugin_logic_bus_toAxi4_aw_valid = LsuL1Plugin_logic_bus_toAxi4_awFiltred_rValid;
  assign LsuL1Plugin_logic_bus_toAxi4_aw_payload_last = LsuL1Plugin_logic_bus_toAxi4_awFiltred_rData_last;
  assign LsuL1Plugin_logic_bus_toAxi4_aw_payload_fragment_address = LsuL1Plugin_logic_bus_toAxi4_awFiltred_rData_fragment_address;
  assign LsuL1Plugin_logic_bus_toAxi4_aw_payload_fragment_data = LsuL1Plugin_logic_bus_toAxi4_awFiltred_rData_fragment_data;
  assign LsuL1Axi4Plugin_logic_axi_aw_valid = LsuL1Plugin_logic_bus_toAxi4_aw_valid;
  assign LsuL1Axi4Plugin_logic_axi_aw_payload_addr = LsuL1Plugin_logic_bus_toAxi4_aw_payload_fragment_address;
  assign LsuL1Axi4Plugin_logic_axi_aw_payload_cache = 4'b1111;
  assign LsuL1Axi4Plugin_logic_axi_aw_payload_prot = 3'b010;
  assign LsuL1Axi4Plugin_logic_axi_aw_payload_len = 8'h07;
  assign LsuL1Axi4Plugin_logic_axi_aw_payload_size = 3'b011;
  assign LsuL1Axi4Plugin_logic_axi_aw_payload_burst = 2'b01;
  assign LsuL1Plugin_logic_bus_toAxi4_aw_ready = LsuL1Axi4Plugin_logic_axi_aw_ready;
  assign _zz_LsuL1Plugin_logic_bus_toAxi4_wRaw_ready = (! LsuL1Plugin_logic_bus_toAxi4_awFiltred_valid);
  assign LsuL1Plugin_logic_bus_toAxi4_w_valid = (LsuL1Plugin_logic_bus_toAxi4_wRaw_valid && _zz_LsuL1Plugin_logic_bus_toAxi4_wRaw_ready);
  assign LsuL1Plugin_logic_bus_toAxi4_wRaw_ready = (LsuL1Plugin_logic_bus_toAxi4_w_ready && _zz_LsuL1Plugin_logic_bus_toAxi4_wRaw_ready);
  assign LsuL1Plugin_logic_bus_toAxi4_w_payload_last = LsuL1Plugin_logic_bus_toAxi4_wRaw_payload_last;
  assign LsuL1Plugin_logic_bus_toAxi4_w_payload_fragment_address = LsuL1Plugin_logic_bus_toAxi4_wRaw_payload_fragment_address;
  assign LsuL1Plugin_logic_bus_toAxi4_w_payload_fragment_data = LsuL1Plugin_logic_bus_toAxi4_wRaw_payload_fragment_data;
  assign LsuL1Axi4Plugin_logic_axi_w_valid = LsuL1Plugin_logic_bus_toAxi4_w_valid;
  assign LsuL1Axi4Plugin_logic_axi_w_payload_data = LsuL1Plugin_logic_bus_toAxi4_w_payload_fragment_data;
  assign LsuL1Axi4Plugin_logic_axi_w_payload_strb = 8'hff;
  assign LsuL1Axi4Plugin_logic_axi_w_payload_last = LsuL1Plugin_logic_bus_toAxi4_w_payload_last;
  assign LsuL1Plugin_logic_bus_toAxi4_w_ready = LsuL1Axi4Plugin_logic_axi_w_ready;
  assign LsuL1Plugin_logic_bus_write_rsp_valid = LsuL1Axi4Plugin_logic_axi_b_valid;
  assign LsuL1Plugin_logic_bus_write_rsp_payload_error = (! (LsuL1Axi4Plugin_logic_axi_b_payload_resp == 2'b00));
  assign LsuL1Axi4Plugin_logic_axi_b_ready = 1'b1;
  always @(*) begin
    CsrAccessPlugin_bus_decode_exception = 1'b0;
    if(when_PrivilegedPlugin_l887) begin
      CsrAccessPlugin_bus_decode_exception = 1'b1;
    end
    if(when_CsrAccessPlugin_l157) begin
      if(when_MmuPlugin_l223) begin
        CsrAccessPlugin_bus_decode_exception = 1'b1;
      end
    end
    if(when_CsrAccessPlugin_l157_2) begin
      if(when_CsrService_l121) begin
        CsrAccessPlugin_bus_decode_exception = 1'b1;
      end
    end
    if(when_CsrAccessPlugin_l157_3) begin
      if(when_CsrService_l121_1) begin
        CsrAccessPlugin_bus_decode_exception = 1'b1;
      end
    end
    if(when_CsrAccessPlugin_l157_4) begin
      if(when_CsrService_l121_2) begin
        CsrAccessPlugin_bus_decode_exception = 1'b1;
      end
    end
    if(when_CsrAccessPlugin_l157_5) begin
      if(when_CsrService_l121_3) begin
        CsrAccessPlugin_bus_decode_exception = 1'b1;
      end
    end
    if(when_CsrAccessPlugin_l157_6) begin
      if(when_CsrService_l198) begin
        if(when_CsrService_l199) begin
          CsrAccessPlugin_bus_decode_exception = 1'b1;
        end
      end
    end
    if(when_CsrAccessPlugin_l157_7) begin
      if(when_CsrService_l121_4) begin
        CsrAccessPlugin_bus_decode_exception = 1'b1;
      end
    end
    if(when_CsrAccessPlugin_l157_8) begin
      if(when_CsrService_l121_5) begin
        CsrAccessPlugin_bus_decode_exception = 1'b1;
      end
    end
    if(when_CsrAccessPlugin_l157_9) begin
      if(when_PerformanceCounterPlugin_l327) begin
        if(when_PerformanceCounterPlugin_l328) begin
          CsrAccessPlugin_bus_decode_exception = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    CsrAccessPlugin_bus_decode_trap = 1'b0;
    if(when_CsrAccessPlugin_l157) begin
      if(!when_MmuPlugin_l223) begin
        CsrAccessPlugin_bus_decode_trap = 1'b1;
      end
    end
    if(when_CsrAccessPlugin_l157_1) begin
      if(CsrAccessPlugin_bus_decode_write) begin
        CsrAccessPlugin_bus_decode_trap = 1'b1;
      end
    end
    if(when_CsrAccessPlugin_l157_10) begin
      if(CsrAccessPlugin_bus_decode_write) begin
        CsrAccessPlugin_bus_decode_trap = 1'b1;
      end
    end
  end

  always @(*) begin
    CsrAccessPlugin_bus_decode_trapCode = 4'bxxxx;
    if(when_CsrAccessPlugin_l157) begin
      if(!when_MmuPlugin_l223) begin
        CsrAccessPlugin_bus_decode_trapCode = 4'b0110;
      end
    end
    if(when_CsrAccessPlugin_l157_1) begin
      if(CsrAccessPlugin_bus_decode_write) begin
        CsrAccessPlugin_bus_decode_trapCode = 4'b0101;
      end
    end
    if(when_CsrAccessPlugin_l157_10) begin
      if(CsrAccessPlugin_bus_decode_write) begin
        CsrAccessPlugin_bus_decode_trapCode = 4'b0101;
      end
    end
  end

  assign CsrAccessPlugin_bus_decode_fence = 1'b0;
  always @(*) begin
    CsrAccessPlugin_bus_read_halt = 1'b0;
    if(when_CsrRamPlugin_l90) begin
      CsrAccessPlugin_bus_read_halt = 1'b1;
    end
  end

  always @(*) begin
    CsrAccessPlugin_bus_write_halt = 1'b0;
    if(when_CsrRamPlugin_l101) begin
      CsrAccessPlugin_bus_write_halt = 1'b1;
    end
    if(when_CsrAccessPlugin_l349_3) begin
      if(when_PerformanceCounterPlugin_l357) begin
        if(when_PerformanceCounterPlugin_l359) begin
          CsrAccessPlugin_bus_write_halt = 1'b1;
        end
      end
    end
  end

  assign FetchL1Plugin_logic_banks_0_read_rsp = FetchL1Plugin_logic_banks_0_mem_spinal_port1;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_WORDS_0 = FetchL1Plugin_logic_banks_0_read_rsp;
  assign FetchL1Plugin_logic_banks_1_read_rsp = FetchL1Plugin_logic_banks_1_mem_spinal_port1;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_WORDS_1 = FetchL1Plugin_logic_banks_1_read_rsp;
  always @(*) begin
    FetchL1Plugin_logic_waysWrite_mask = 2'b00;
    if(when_FetchL1Plugin_l204) begin
      FetchL1Plugin_logic_waysWrite_mask = 2'b11;
    end
    if(FetchL1Plugin_logic_invalidate_done) begin
      if(when_FetchL1Plugin_l304) begin
        FetchL1Plugin_logic_waysWrite_mask[FetchL1Plugin_logic_refill_onRsp_wayToAllocate] = 1'b1;
      end
    end
  end

  always @(*) begin
    FetchL1Plugin_logic_waysWrite_address = 6'bxxxxxx;
    if(when_FetchL1Plugin_l204) begin
      FetchL1Plugin_logic_waysWrite_address = FetchL1Plugin_logic_invalidate_counter[5:0];
    end
    if(FetchL1Plugin_logic_invalidate_done) begin
      FetchL1Plugin_logic_waysWrite_address = FetchL1Plugin_logic_refill_onRsp_address[11 : 6];
    end
  end

  always @(*) begin
    FetchL1Plugin_logic_waysWrite_tag_loaded = 1'bx;
    if(when_FetchL1Plugin_l204) begin
      FetchL1Plugin_logic_waysWrite_tag_loaded = 1'b0;
    end
    if(FetchL1Plugin_logic_invalidate_done) begin
      FetchL1Plugin_logic_waysWrite_tag_loaded = 1'b1;
    end
  end

  always @(*) begin
    FetchL1Plugin_logic_waysWrite_tag_error = 1'bx;
    if(FetchL1Plugin_logic_invalidate_done) begin
      FetchL1Plugin_logic_waysWrite_tag_error = (FetchL1Plugin_logic_bus_rsp_valid && FetchL1Plugin_logic_bus_rsp_payload_error);
    end
  end

  always @(*) begin
    FetchL1Plugin_logic_waysWrite_tag_address = 20'bxxxxxxxxxxxxxxxxxxxx;
    if(FetchL1Plugin_logic_invalidate_done) begin
      FetchL1Plugin_logic_waysWrite_tag_address = FetchL1Plugin_logic_refill_onRsp_address[31 : 12];
    end
  end

  assign _zz_FetchL1Plugin_logic_ways_0_read_rsp_loaded = FetchL1Plugin_logic_ways_0_mem_spinal_port1;
  assign FetchL1Plugin_logic_ways_0_read_rsp_loaded = _zz_FetchL1Plugin_logic_ways_0_read_rsp_loaded[0];
  assign FetchL1Plugin_logic_ways_0_read_rsp_error = _zz_FetchL1Plugin_logic_ways_0_read_rsp_loaded[1];
  assign FetchL1Plugin_logic_ways_0_read_rsp_address = _zz_FetchL1Plugin_logic_ways_0_read_rsp_loaded[21 : 2];
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_loaded = FetchL1Plugin_logic_ways_0_read_rsp_loaded;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_error = FetchL1Plugin_logic_ways_0_read_rsp_error;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_address = FetchL1Plugin_logic_ways_0_read_rsp_address;
  assign _zz_FetchL1Plugin_logic_ways_1_read_rsp_loaded = FetchL1Plugin_logic_ways_1_mem_spinal_port1;
  assign FetchL1Plugin_logic_ways_1_read_rsp_loaded = _zz_FetchL1Plugin_logic_ways_1_read_rsp_loaded[0];
  assign FetchL1Plugin_logic_ways_1_read_rsp_error = _zz_FetchL1Plugin_logic_ways_1_read_rsp_loaded[1];
  assign FetchL1Plugin_logic_ways_1_read_rsp_address = _zz_FetchL1Plugin_logic_ways_1_read_rsp_loaded[21 : 2];
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_loaded = FetchL1Plugin_logic_ways_1_read_rsp_loaded;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_error = FetchL1Plugin_logic_ways_1_read_rsp_error;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_address = FetchL1Plugin_logic_ways_1_read_rsp_address;
  assign FetchL1Plugin_logic_plru_read_rsp_0 = FetchL1Plugin_logic_plru_mem_spinal_port1[0 : 0];
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_PLRU_READ_0 = FetchL1Plugin_logic_plru_read_rsp_0;
  assign FetchL1Plugin_logic_invalidate_cmd_valid = (|TrapPlugin_logic_fetchL1Invalidate_0_cmd_valid);
  always @(*) begin
    FetchL1Plugin_logic_invalidate_canStart = 1'b1;
    if(when_FetchL1Plugin_l268) begin
      FetchL1Plugin_logic_invalidate_canStart = 1'b0;
    end
  end

  assign FetchL1Plugin_logic_invalidate_counterIncr = (FetchL1Plugin_logic_invalidate_counter + 7'h01);
  assign FetchL1Plugin_logic_invalidate_done = FetchL1Plugin_logic_invalidate_counter[6];
  assign FetchL1Plugin_logic_invalidate_last = FetchL1Plugin_logic_invalidate_counterIncr[6];
  assign when_FetchL1Plugin_l204 = (! FetchL1Plugin_logic_invalidate_done);
  assign when_FetchL1Plugin_l211 = ((FetchL1Plugin_logic_invalidate_done && FetchL1Plugin_logic_invalidate_cmd_valid) && FetchL1Plugin_logic_invalidate_canStart);
  always @(*) begin
    TrapPlugin_logic_fetchL1Invalidate_0_cmd_ready = 1'b0;
    if(when_FetchL1Plugin_l216) begin
      if(FetchL1Plugin_logic_invalidate_last) begin
        TrapPlugin_logic_fetchL1Invalidate_0_cmd_ready = 1'b1;
      end
    end
  end

  assign when_FetchL1Plugin_l216 = (! FetchL1Plugin_logic_invalidate_done);
  assign fetch_logic_ctrls_0_haltRequest_FetchL1Plugin_l217 = _zz_fetch_logic_ctrls_0_haltRequest_FetchL1Plugin_l217;
  assign FetchL1Plugin_logic_refill_slots_0_askCmd = (FetchL1Plugin_logic_refill_slots_0_valid && (! FetchL1Plugin_logic_refill_slots_0_cmdSent));
  assign FetchL1Plugin_logic_refill_hazard = (|(FetchL1Plugin_logic_refill_slots_0_valid && (FetchL1Plugin_logic_refill_slots_0_address[11 : 6] == FetchL1Plugin_logic_refill_start_address[11 : 6])));
  assign when_FetchL1Plugin_l255 = ((FetchL1Plugin_logic_refill_start_valid && FetchL1Plugin_logic_invalidate_done) && (! FetchL1Plugin_logic_refill_hazard));
  assign when_FetchL1Plugin_l268 = ((|FetchL1Plugin_logic_refill_slots_0_valid) || FetchL1Plugin_logic_refill_start_valid);
  assign FetchL1Plugin_logic_refill_onCmd_propoedOh = (FetchL1Plugin_logic_refill_slots_0_askCmd && 1'b1);
  assign when_FetchL1Plugin_l276 = (! FetchL1Plugin_logic_refill_onCmd_locked);
  assign FetchL1Plugin_logic_refill_onCmd_oh = (FetchL1Plugin_logic_refill_onCmd_locked ? FetchL1Plugin_logic_refill_onCmd_lockedOh : FetchL1Plugin_logic_refill_onCmd_propoedOh);
  assign FetchL1Plugin_logic_bus_cmd_valid = (|FetchL1Plugin_logic_refill_onCmd_oh);
  assign FetchL1Plugin_logic_bus_cmd_payload_address = {FetchL1Plugin_logic_refill_slots_0_address[31 : 6],6'h0};
  assign FetchL1Plugin_logic_bus_cmd_payload_io = FetchL1Plugin_logic_refill_slots_0_isIo;
  assign FetchL1Plugin_logic_refill_onRsp_holdHarts = ((|FetchL1Plugin_logic_waysWrite_mask) || (|((FetchL1Plugin_logic_refill_slots_0_valid && (FetchL1Plugin_logic_refill_slots_0_address[11 : 6] == fetch_logic_ctrls_0_down_Fetch_WORD_PC[11 : 6])) && (! (1'b1 && (fetch_logic_ctrls_0_down_Fetch_WORD_PC[5 : 3] < FetchL1Plugin_logic_refill_onRsp_wordIndex))))));
  assign fetch_logic_ctrls_0_haltRequest_FetchL1Plugin_l297 = FetchL1Plugin_logic_refill_onRsp_holdHarts;
  assign FetchL1Plugin_logic_bus_rsp_fire = (FetchL1Plugin_logic_bus_rsp_valid && FetchL1Plugin_logic_bus_rsp_ready);
  assign FetchL1Plugin_logic_refill_onRsp_wayToAllocate = FetchL1Plugin_logic_refill_slots_0_wayToAllocate;
  assign FetchL1Plugin_logic_refill_onRsp_address = FetchL1Plugin_logic_refill_slots_0_address;
  assign when_FetchL1Plugin_l304 = (FetchL1Plugin_logic_bus_rsp_valid && (FetchL1Plugin_logic_refill_onRsp_firstCycle || FetchL1Plugin_logic_bus_rsp_payload_error));
  assign FetchL1Plugin_logic_banks_0_write_valid = (FetchL1Plugin_logic_bus_rsp_valid && (FetchL1Plugin_logic_refill_onRsp_wayToAllocate == 1'b0));
  assign FetchL1Plugin_logic_banks_0_write_payload_address = {FetchL1Plugin_logic_refill_onRsp_address[11 : 6],FetchL1Plugin_logic_refill_onRsp_wordIndex};
  assign FetchL1Plugin_logic_banks_0_write_payload_data = FetchL1Plugin_logic_bus_rsp_payload_data;
  assign FetchL1Plugin_logic_banks_1_write_valid = (FetchL1Plugin_logic_bus_rsp_valid && (FetchL1Plugin_logic_refill_onRsp_wayToAllocate == 1'b1));
  assign FetchL1Plugin_logic_banks_1_write_payload_address = {FetchL1Plugin_logic_refill_onRsp_address[11 : 6],FetchL1Plugin_logic_refill_onRsp_wordIndex};
  assign FetchL1Plugin_logic_banks_1_write_payload_data = FetchL1Plugin_logic_bus_rsp_payload_data;
  assign FetchL1Plugin_logic_bus_rsp_ready = 1'b1;
  assign when_FetchL1Plugin_l330 = (FetchL1Plugin_logic_refill_onRsp_wordIndex == 3'b111);
  assign FetchL1Plugin_logic_cmd_doIt = (fetch_logic_ctrls_1_up_ready || ((! fetch_logic_ctrls_1_up_valid) && 1'b1));
  assign FetchL1Plugin_logic_banks_0_read_cmd_valid = FetchL1Plugin_logic_cmd_doIt;
  assign FetchL1Plugin_logic_banks_0_read_cmd_payload = fetch_logic_ctrls_0_down_Fetch_WORD_PC[11 : 3];
  assign FetchL1Plugin_logic_banks_1_read_cmd_valid = FetchL1Plugin_logic_cmd_doIt;
  assign FetchL1Plugin_logic_banks_1_read_cmd_payload = fetch_logic_ctrls_0_down_Fetch_WORD_PC[11 : 3];
  assign FetchL1Plugin_logic_ways_0_read_cmd_valid = FetchL1Plugin_logic_cmd_doIt;
  assign FetchL1Plugin_logic_ways_0_read_cmd_payload = fetch_logic_ctrls_0_down_Fetch_WORD_PC[11 : 6];
  assign FetchL1Plugin_logic_ways_1_read_cmd_valid = FetchL1Plugin_logic_cmd_doIt;
  assign FetchL1Plugin_logic_ways_1_read_cmd_payload = fetch_logic_ctrls_0_down_Fetch_WORD_PC[11 : 6];
  assign FetchL1Plugin_logic_plru_read_cmd_valid = FetchL1Plugin_logic_cmd_doIt;
  assign FetchL1Plugin_logic_plru_read_cmd_payload = fetch_logic_ctrls_0_down_Fetch_WORD_PC[11 : 6];
  assign fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_VALID = (FetchL1Plugin_logic_plru_write_valid && (FetchL1Plugin_logic_plru_write_payload_address == FetchL1Plugin_logic_plru_read_cmd_payload));
  assign fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_0 = FetchL1Plugin_logic_plru_write_payload_data_0;
  assign fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE = (|FetchL1Plugin_logic_waysWrite_mask);
  assign fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE_ADDRESS = FetchL1Plugin_logic_waysWrite_address;
  always @(*) begin
    fetch_logic_ctrls_1_down_FetchL1Plugin_logic_PLRU_BYPASSED_0 = fetch_logic_ctrls_1_down_FetchL1Plugin_logic_PLRU_READ_0;
    if(fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_VALID) begin
      fetch_logic_ctrls_1_down_FetchL1Plugin_logic_PLRU_BYPASSED_0 = fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_0;
    end
  end

  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_0 = _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_0;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_1 = _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_1;
  assign fetch_logic_ctrls_2_down_Fetch_WORD = ((fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_0 ? fetch_logic_ctrls_2_down_FetchL1Plugin_logic_BANKS_MUXES_0 : 32'h0) | (fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_1 ? fetch_logic_ctrls_2_down_FetchL1Plugin_logic_BANKS_MUXES_1 : 32'h0));
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_HAZARD = (fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE && (fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE_ADDRESS == fetch_logic_ctrls_1_down_Fetch_WORD_PC[11 : 6]));
  assign FetchL1Plugin_logic_hits_w_0_indirect_wayTlbHits_0 = ((fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_address == fetch_logic_ctrls_1_down_MMU_WAYS_PHYSICAL_0[31 : 12]) && fetch_logic_ctrls_1_down_MMU_WAYS_OH[0]);
  assign FetchL1Plugin_logic_hits_w_0_indirect_wayTlbHits_1 = ((fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_address == fetch_logic_ctrls_1_down_MMU_WAYS_PHYSICAL_1[31 : 12]) && fetch_logic_ctrls_1_down_MMU_WAYS_OH[1]);
  assign FetchL1Plugin_logic_hits_w_0_indirect_wayTlbHits_2 = ((fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_address == fetch_logic_ctrls_1_down_MMU_WAYS_PHYSICAL_2[31 : 12]) && fetch_logic_ctrls_1_down_MMU_WAYS_OH[2]);
  assign FetchL1Plugin_logic_hits_w_0_indirect_translatedHits = (|{FetchL1Plugin_logic_hits_w_0_indirect_wayTlbHits_2,{FetchL1Plugin_logic_hits_w_0_indirect_wayTlbHits_1,FetchL1Plugin_logic_hits_w_0_indirect_wayTlbHits_0}});
  assign FetchL1Plugin_logic_hits_w_0_indirect_bypassHits = (_zz_FetchL1Plugin_logic_hits_w_0_indirect_bypassHits == _zz_FetchL1Plugin_logic_hits_w_0_indirect_bypassHits_1);
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HITS_0 = ((fetch_logic_ctrls_1_down_MMU_BYPASS_TRANSLATION ? FetchL1Plugin_logic_hits_w_0_indirect_bypassHits : FetchL1Plugin_logic_hits_w_0_indirect_translatedHits) && fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_loaded);
  assign FetchL1Plugin_logic_hits_w_1_indirect_wayTlbHits_0 = ((fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_address == fetch_logic_ctrls_1_down_MMU_WAYS_PHYSICAL_0[31 : 12]) && fetch_logic_ctrls_1_down_MMU_WAYS_OH[0]);
  assign FetchL1Plugin_logic_hits_w_1_indirect_wayTlbHits_1 = ((fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_address == fetch_logic_ctrls_1_down_MMU_WAYS_PHYSICAL_1[31 : 12]) && fetch_logic_ctrls_1_down_MMU_WAYS_OH[1]);
  assign FetchL1Plugin_logic_hits_w_1_indirect_wayTlbHits_2 = ((fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_address == fetch_logic_ctrls_1_down_MMU_WAYS_PHYSICAL_2[31 : 12]) && fetch_logic_ctrls_1_down_MMU_WAYS_OH[2]);
  assign FetchL1Plugin_logic_hits_w_1_indirect_translatedHits = (|{FetchL1Plugin_logic_hits_w_1_indirect_wayTlbHits_2,{FetchL1Plugin_logic_hits_w_1_indirect_wayTlbHits_1,FetchL1Plugin_logic_hits_w_1_indirect_wayTlbHits_0}});
  assign FetchL1Plugin_logic_hits_w_1_indirect_bypassHits = (_zz_FetchL1Plugin_logic_hits_w_1_indirect_bypassHits == _zz_FetchL1Plugin_logic_hits_w_1_indirect_bypassHits_1);
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HITS_1 = ((fetch_logic_ctrls_1_down_MMU_BYPASS_TRANSLATION ? FetchL1Plugin_logic_hits_w_1_indirect_bypassHits : FetchL1Plugin_logic_hits_w_1_indirect_translatedHits) && fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_loaded);
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HIT = (|{fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HITS_1,fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HITS_0});
  assign FetchL1Plugin_logic_ctrl_pmaPort_cmd_address = fetch_logic_ctrls_2_down_MMU_TRANSLATED;
  assign FetchL1Plugin_logic_ctrl_plruLogic_core_evict_logic_0_state = FetchL1Plugin_logic_ctrl_plruLogic_core_io_context_state_0[0];
  assign FetchL1Plugin_logic_ctrl_plruLogic_core_evict_sel_0 = (! FetchL1Plugin_logic_ctrl_plruLogic_core_evict_logic_0_state);
  assign FetchL1Plugin_logic_ctrl_plruLogic_core_io_evict_id = FetchL1Plugin_logic_ctrl_plruLogic_core_evict_sel_0;
  assign FetchL1Plugin_logic_ctrl_plruLogic_core_io_update_state_0[0] = FetchL1Plugin_logic_ctrl_plruLogic_core_io_update_id[0];
  assign FetchL1Plugin_logic_ctrl_plruLogic_core_io_context_state_0 = fetch_logic_ctrls_2_down_FetchL1Plugin_logic_PLRU_BYPASSED_0;
  assign FetchL1Plugin_logic_ctrl_plruLogic_core_io_update_id = fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_1;
  always @(*) begin
    FetchL1Plugin_logic_plru_write_valid = FetchL1Plugin_logic_ctrl_plruLogic_buffer_regNext_valid;
    if(when_FetchL1Plugin_l558) begin
      FetchL1Plugin_logic_plru_write_valid = 1'b1;
    end
  end

  always @(*) begin
    FetchL1Plugin_logic_plru_write_payload_address = FetchL1Plugin_logic_ctrl_plruLogic_buffer_regNext_payload_address;
    if(when_FetchL1Plugin_l558) begin
      FetchL1Plugin_logic_plru_write_payload_address = FetchL1Plugin_logic_invalidate_counter[5:0];
    end
  end

  always @(*) begin
    FetchL1Plugin_logic_plru_write_payload_data_0 = FetchL1Plugin_logic_ctrl_plruLogic_buffer_regNext_payload_data_0;
    if(when_FetchL1Plugin_l558) begin
      FetchL1Plugin_logic_plru_write_payload_data_0 = _zz_FetchL1Plugin_logic_plru_write_payload_data_0[0 : 0];
    end
  end

  assign FetchL1Plugin_logic_ctrl_plruLogic_buffer_valid = (fetch_logic_ctrls_2_up_isValid && fetch_logic_ctrls_2_up_isReady);
  assign FetchL1Plugin_logic_ctrl_plruLogic_buffer_payload_address = fetch_logic_ctrls_2_down_Fetch_WORD_PC[11 : 6];
  assign FetchL1Plugin_logic_ctrl_plruLogic_buffer_payload_data_0 = FetchL1Plugin_logic_ctrl_plruLogic_core_io_update_state_0;
  assign FetchL1Plugin_logic_refill_start_wayToAllocate = FetchL1Plugin_logic_ctrl_plruLogic_core_io_evict_id;
  assign FetchL1Plugin_logic_ctrl_dataAccessFault = (_zz_FetchL1Plugin_logic_ctrl_dataAccessFault[0] && (! fetch_logic_ctrls_2_down_FetchL1Plugin_logic_HAZARD));
  always @(*) begin
    FetchL1Plugin_logic_trapPort_valid = 1'b0;
    if(when_FetchL1Plugin_l474) begin
      FetchL1Plugin_logic_trapPort_valid = 1'b1;
    end
    if(when_FetchL1Plugin_l480) begin
      FetchL1Plugin_logic_trapPort_valid = 1'b1;
    end
    if(when_FetchL1Plugin_l487) begin
      FetchL1Plugin_logic_trapPort_valid = 1'b1;
    end
    if(fetch_logic_ctrls_2_down_MMU_ACCESS_FAULT) begin
      FetchL1Plugin_logic_trapPort_valid = 1'b1;
    end
    if(fetch_logic_ctrls_2_down_MMU_REFILL) begin
      FetchL1Plugin_logic_trapPort_valid = 1'b1;
    end
    if(fetch_logic_ctrls_2_down_MMU_HAZARD) begin
      FetchL1Plugin_logic_trapPort_valid = 1'b1;
    end
    if(fetch_logic_ctrls_2_down_Fetch_PC_FAULT) begin
      FetchL1Plugin_logic_trapPort_valid = 1'b1;
    end
    if(when_FetchL1Plugin_l533) begin
      FetchL1Plugin_logic_trapPort_valid = 1'b0;
    end
  end

  assign FetchL1Plugin_logic_trapPort_payload_tval = fetch_logic_ctrls_2_down_Fetch_WORD_PC;
  always @(*) begin
    FetchL1Plugin_logic_trapPort_payload_exception = 1'bx;
    if(when_FetchL1Plugin_l474) begin
      FetchL1Plugin_logic_trapPort_payload_exception = 1'b0;
    end
    if(when_FetchL1Plugin_l480) begin
      FetchL1Plugin_logic_trapPort_payload_exception = 1'b1;
    end
    if(when_FetchL1Plugin_l487) begin
      FetchL1Plugin_logic_trapPort_payload_exception = 1'b1;
    end
    if(fetch_logic_ctrls_2_down_MMU_ACCESS_FAULT) begin
      FetchL1Plugin_logic_trapPort_payload_exception = 1'b1;
    end
    if(fetch_logic_ctrls_2_down_MMU_REFILL) begin
      FetchL1Plugin_logic_trapPort_payload_exception = 1'b0;
    end
    if(fetch_logic_ctrls_2_down_MMU_HAZARD) begin
      FetchL1Plugin_logic_trapPort_payload_exception = 1'b0;
    end
    if(fetch_logic_ctrls_2_down_Fetch_PC_FAULT) begin
      FetchL1Plugin_logic_trapPort_payload_exception = 1'b1;
    end
  end

  always @(*) begin
    FetchL1Plugin_logic_trapPort_payload_code = 4'bxxxx;
    if(when_FetchL1Plugin_l474) begin
      FetchL1Plugin_logic_trapPort_payload_code = 4'b0100;
    end
    if(when_FetchL1Plugin_l480) begin
      FetchL1Plugin_logic_trapPort_payload_code = 4'b0001;
    end
    if(when_FetchL1Plugin_l487) begin
      FetchL1Plugin_logic_trapPort_payload_code = 4'b1100;
    end
    if(fetch_logic_ctrls_2_down_MMU_ACCESS_FAULT) begin
      FetchL1Plugin_logic_trapPort_payload_code = 4'b0001;
    end
    if(fetch_logic_ctrls_2_down_MMU_REFILL) begin
      FetchL1Plugin_logic_trapPort_payload_code = 4'b0111;
    end
    if(fetch_logic_ctrls_2_down_MMU_HAZARD) begin
      FetchL1Plugin_logic_trapPort_payload_code = 4'b0100;
    end
    if(fetch_logic_ctrls_2_down_Fetch_PC_FAULT) begin
      FetchL1Plugin_logic_trapPort_payload_code = 4'b0001;
      if(when_FetchL1Plugin_l520) begin
        FetchL1Plugin_logic_trapPort_payload_code = 4'b1100;
      end
    end
  end

  assign _zz_60 = zz_FetchL1Plugin_logic_trapPort_payload_arg(1'b0);
  always @(*) FetchL1Plugin_logic_trapPort_payload_arg = _zz_60;
  always @(*) begin
    FetchL1Plugin_logic_ctrl_allowRefill = ((! fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HIT) && (! fetch_logic_ctrls_2_down_FetchL1Plugin_logic_HAZARD));
    if(when_FetchL1Plugin_l480) begin
      FetchL1Plugin_logic_ctrl_allowRefill = 1'b0;
    end
    if(when_FetchL1Plugin_l487) begin
      FetchL1Plugin_logic_ctrl_allowRefill = 1'b0;
    end
    if(fetch_logic_ctrls_2_down_MMU_ACCESS_FAULT) begin
      FetchL1Plugin_logic_ctrl_allowRefill = 1'b0;
    end
    if(fetch_logic_ctrls_2_down_MMU_REFILL) begin
      FetchL1Plugin_logic_ctrl_allowRefill = 1'b0;
    end
    if(fetch_logic_ctrls_2_down_MMU_HAZARD) begin
      FetchL1Plugin_logic_ctrl_allowRefill = 1'b0;
    end
    if(fetch_logic_ctrls_2_down_Fetch_PC_FAULT) begin
      FetchL1Plugin_logic_ctrl_allowRefill = 1'b0;
    end
  end

  assign when_FetchL1Plugin_l474 = ((! fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HIT) || fetch_logic_ctrls_2_down_FetchL1Plugin_logic_HAZARD);
  assign when_FetchL1Plugin_l480 = ((FetchL1Plugin_logic_ctrl_dataAccessFault || FetchL1Plugin_logic_ctrl_pmaPort_rsp_fault) || fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_ACCESS_FAULT);
  assign when_FetchL1Plugin_l487 = (fetch_logic_ctrls_2_down_MMU_PAGE_FAULT || (! fetch_logic_ctrls_2_down_MMU_ALLOW_EXECUTE));
  assign when_FetchL1Plugin_l520 = (! fetch_logic_ctrls_2_down_MMU_BYPASS_TRANSLATION);
  always @(*) begin
    FetchL1Plugin_logic_refill_start_valid = (FetchL1Plugin_logic_ctrl_allowRefill && (! FetchL1Plugin_logic_ctrl_trapSent));
    if(when_FetchL1Plugin_l537) begin
      FetchL1Plugin_logic_refill_start_valid = 1'b0;
    end
  end

  assign FetchL1Plugin_logic_refill_start_address = fetch_logic_ctrls_2_down_MMU_TRANSLATED;
  assign FetchL1Plugin_logic_refill_start_isIo = FetchL1Plugin_logic_ctrl_pmaPort_rsp_io;
  assign fetch_logic_ctrls_2_down_TRAP = (FetchL1Plugin_logic_trapPort_valid || FetchL1Plugin_logic_ctrl_trapSent);
  assign when_FetchL1Plugin_l533 = ((! fetch_logic_ctrls_2_up_isValid) || FetchL1Plugin_logic_ctrl_trapSent);
  assign when_FetchL1Plugin_l537 = ((! fetch_logic_ctrls_2_up_isValid) && 1'b1);
  assign when_FetchL1Plugin_l541 = (((! fetch_logic_ctrls_2_up_isValid) || fetch_logic_ctrls_2_down_isReady) || fetch_logic_ctrls_2_up_isCanceling);
  assign when_FetchL1Plugin_l549 = (fetch_logic_ctrls_2_up_isValid && (! fetch_logic_ctrls_2_down_TRAP));
  assign FetchL1Plugin_logic_events_access = fetch_logic_ctrls_2_up_isMoving;
  assign FetchL1Plugin_logic_events_miss = (fetch_logic_ctrls_2_up_isMoving && FetchL1Plugin_logic_ctrl_allowRefill);
  assign FetchL1Plugin_logic_events_waiting = FetchL1Plugin_logic_ctrl_onEvents_waiting;
  assign when_FetchL1Plugin_l558 = (! FetchL1Plugin_logic_invalidate_done);
  assign LsuPlugin_logic_frontend_defaultsDecodings_0 = 1'b0;
  assign LsuPlugin_logic_frontend_defaultsDecodings_1 = 1'b0;
  assign LsuPlugin_logic_frontend_defaultsDecodings_2 = 1'b0;
  assign LsuPlugin_logic_frontend_defaultsDecodings_3 = 1'b0;
  assign LsuPlugin_logic_frontend_defaultsDecodings_4 = 1'b0;
  assign LsuPlugin_logic_frontend_defaultsDecodings_5 = 1'b0;
  always @(*) begin
    LsuPlugin_logic_cbmCsr_invalIntoClean = 1'b0;
    if(when_LsuPlugin_l226) begin
      LsuPlugin_logic_cbmCsr_invalIntoClean = 1'b1;
    end
    if(when_LsuPlugin_l226_1) begin
      LsuPlugin_logic_cbmCsr_invalIntoClean = 1'b1;
    end
  end

  always @(*) begin
    PrivilegedPlugin_logic_harts_0_xretAwayFromMachine = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_WAIT : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
        if(when_TrapPlugin_l712) begin
          PrivilegedPlugin_logic_harts_0_xretAwayFromMachine = 1'b1;
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    PrivilegedPlugin_logic_harts_0_int_pending = 1'b0;
    if(TrapPlugin_logic_harts_0_interrupt_pendingInterrupt) begin
      PrivilegedPlugin_logic_harts_0_int_pending = 1'b1;
    end
  end

  assign PrivilegedPlugin_logic_harts_0_withMachinePrivilege = (2'b11 <= PrivilegedPlugin_logic_harts_0_privilege);
  assign PrivilegedPlugin_logic_harts_0_withSupervisorPrivilege = (2'b01 <= PrivilegedPlugin_logic_harts_0_privilege);
  assign PrivilegedPlugin_logic_harts_0_hartRunning = 1'b1;
  assign PrivilegedPlugin_logic_harts_0_debugMode = (! PrivilegedPlugin_logic_harts_0_hartRunning);
  always @(*) begin
    PrivilegedPlugin_logic_harts_0_m_status_sd = 1'b0;
    if(when_PrivilegedPlugin_l573) begin
      PrivilegedPlugin_logic_harts_0_m_status_sd = 1'b1;
    end
  end

  assign when_PrivilegedPlugin_l573 = (PrivilegedPlugin_logic_harts_0_m_status_fs == 2'b11);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_12 = (when_CsrService_l232 && _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_13 = (when_CsrService_l232 && REG_CSR_834);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_15 = (when_CsrService_l232 && _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_14);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_17 = (when_CsrService_l232 && _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_16);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_18 = (when_CsrService_l232 && REG_CSR_770);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_20 = (when_CsrService_l232 && _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_19);
  assign _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_0_valid = (PrivilegedPlugin_logic_harts_0_m_ip_mtip && PrivilegedPlugin_logic_harts_0_m_ie_mtie);
  assign _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_1_valid = (PrivilegedPlugin_logic_harts_0_m_ip_msip && PrivilegedPlugin_logic_harts_0_m_ie_msie);
  assign _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_2_valid = (PrivilegedPlugin_logic_harts_0_m_ip_meip && PrivilegedPlugin_logic_harts_0_m_ie_meie);
  always @(*) begin
    PrivilegedPlugin_logic_harts_0_m_topi_interrupt = 4'bxxxx;
    PrivilegedPlugin_logic_harts_0_m_topi_interrupt = TrapPlugin_logic_harts_0_interrupt_xtopi_1_int;
  end

  assign PrivilegedPlugin_logic_harts_0_m_topi_priority = ((PrivilegedPlugin_logic_harts_0_m_topi_interrupt == 4'b0000) ? 1'b0 : 1'b1);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_21 = (when_CsrService_l232 && REG_CSR_4016);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_23 = (when_CsrService_l232 && REG_CSR_322);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_24 = (when_CsrService_l232 && _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_1);
  assign PrivilegedPlugin_logic_harts_0_s_sstc_envcfg_allowUpdate = 1'b0;
  assign PrivilegedPlugin_logic_harts_0_s_sstc_interrupt = 1'b0;
  assign PrivilegedPlugin_logic_harts_0_s_ip_seipOr = (PrivilegedPlugin_logic_harts_0_s_ip_seipSoft || PrivilegedPlugin_logic_harts_0_s_ip_seipInput);
  assign PrivilegedPlugin_logic_harts_0_s_ip_stipOr = (PrivilegedPlugin_logic_harts_0_s_sstc_envcfg_enable ? PrivilegedPlugin_logic_harts_0_s_sstc_interrupt : PrivilegedPlugin_logic_harts_0_s_ip_stipSoft);
  assign PrivilegedPlugin_logic_harts_0_s_ip_seipMasked = (PrivilegedPlugin_logic_harts_0_s_ip_seipOr && PrivilegedPlugin_logic_harts_0_m_ideleg_se);
  assign PrivilegedPlugin_logic_harts_0_s_ip_stipMasked = (PrivilegedPlugin_logic_harts_0_s_ip_stipOr && PrivilegedPlugin_logic_harts_0_m_ideleg_st);
  assign PrivilegedPlugin_logic_harts_0_s_ip_ssipMasked = (PrivilegedPlugin_logic_harts_0_s_ip_ssip && PrivilegedPlugin_logic_harts_0_m_ideleg_ss);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_26 = (when_CsrService_l232 && REG_CSR_260);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_27 = (when_CsrService_l232 && REG_CSR_324);
  assign when_CsrService_l225 = (! PrivilegedPlugin_logic_harts_0_s_sstc_envcfg_enable);
  assign _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_0_valid = (PrivilegedPlugin_logic_harts_0_s_ip_ssip && PrivilegedPlugin_logic_harts_0_s_ie_ssie);
  assign _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_1_valid = (PrivilegedPlugin_logic_harts_0_s_ip_stipOr && PrivilegedPlugin_logic_harts_0_s_ie_stie);
  assign _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_2_valid = (PrivilegedPlugin_logic_harts_0_s_ip_seipOr && PrivilegedPlugin_logic_harts_0_s_ie_seie);
  always @(*) begin
    PrivilegedPlugin_logic_harts_0_s_topi_interrupt = 4'bxxxx;
    PrivilegedPlugin_logic_harts_0_s_topi_interrupt = TrapPlugin_logic_harts_0_interrupt_xtopi_0_int;
  end

  assign PrivilegedPlugin_logic_harts_0_s_topi_priority = ((PrivilegedPlugin_logic_harts_0_s_topi_interrupt == 4'b0000) ? 1'b0 : 1'b1);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_28 = (when_CsrService_l232 && REG_CSR_3504);
  assign PrivilegedPlugin_logic_harts_0_time_accessable = (PrivilegedPlugin_logic_harts_0_withMachinePrivilege || PrivilegedPlugin_logic_harts_0_mcounteren_tm);
  assign PrivilegedPlugin_logic_defaultTrap_csrPrivilege = CsrAccessPlugin_bus_decode_address[9 : 8];
  assign PrivilegedPlugin_logic_defaultTrap_csrReadOnly = (CsrAccessPlugin_bus_decode_address[11 : 10] == 2'b11);
  assign when_PrivilegedPlugin_l887 = ((PrivilegedPlugin_logic_defaultTrap_csrReadOnly && CsrAccessPlugin_bus_decode_write) || (PrivilegedPlugin_logic_harts_0_privilege < PrivilegedPlugin_logic_defaultTrap_csrPrivilege));
  assign GSharePlugin_logic_mem_writes_0_valid = (GSharePlugin_logic_mem_write_valid && 1'b1);
  assign GSharePlugin_logic_mem_writes_0_payload_address = GSharePlugin_logic_mem_write_payload_address;
  assign GSharePlugin_logic_mem_writes_0_payload_data_0 = GSharePlugin_logic_mem_write_payload_data_0;
  assign GSharePlugin_logic_mem_writes_0_payload_data_1 = GSharePlugin_logic_mem_write_payload_data_1;
  assign _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH = fetch_logic_ctrls_0_down_Fetch_WORD_PC[14 : 2];
  assign fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH = ({_zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH[0],{_zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH[1],{_zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH[2],{_zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH[3],{_zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH[4],{_zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH[5],{_zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_1,{_zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_2,_zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_3}}}}}}}} ^ _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_4);
  assign fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_valid = GSharePlugin_logic_mem_write_valid;
  assign fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_address = GSharePlugin_logic_mem_write_payload_address;
  assign fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_data_0 = GSharePlugin_logic_mem_write_payload_data_0;
  assign fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_data_1 = GSharePlugin_logic_mem_write_payload_data_1;
  assign _zz_GSharePlugin_logic_readRsp_readed_0_0 = fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH;
  assign _zz_GSharePlugin_logic_readRsp_readed_0_0_1 = GSharePlugin_logic_mem_banks_0_spinal_port1;
  assign GSharePlugin_logic_readRsp_readed_0_0 = _zz_GSharePlugin_logic_readRsp_readed_0_0_1[1 : 0];
  assign GSharePlugin_logic_readRsp_readed_0_1 = _zz_GSharePlugin_logic_readRsp_readed_0_0_1[3 : 2];
  always @(*) begin
    fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0 = GSharePlugin_logic_readRsp_readed_0_0;
    if(when_GSharePlugin_l100) begin
      fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0 = fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_data_0;
    end
  end

  always @(*) begin
    fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_1 = GSharePlugin_logic_readRsp_readed_0_1;
    if(when_GSharePlugin_l100) begin
      fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_1 = fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_data_1;
    end
  end

  assign when_GSharePlugin_l100 = (fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_valid && (fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_address == fetch_logic_ctrls_1_down_GSharePlugin_logic_HASH));
  always @(*) begin
    BtbPlugin_logic_ras_ptr_pushIt = 1'b0;
    if(BtbPlugin_logic_applyIt_rasLogic_pushValid) begin
      BtbPlugin_logic_ras_ptr_pushIt = 1'b1;
    end
  end

  always @(*) begin
    BtbPlugin_logic_ras_ptr_popIt = 1'b0;
    if(when_BtbPlugin_l246) begin
      BtbPlugin_logic_ras_ptr_popIt = 1'b1;
    end
  end

  assign BtbPlugin_logic_ras_write_valid = BtbPlugin_logic_ras_ptr_pushIt;
  assign BtbPlugin_logic_ras_write_payload_address = BtbPlugin_logic_ras_ptr_push;
  always @(*) begin
    BtbPlugin_logic_ras_write_payload_data = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    BtbPlugin_logic_ras_write_payload_data = (_zz_BtbPlugin_logic_ras_write_payload_data >>> 1'd1);
  end

  assign BtbPlugin_logic_memDp_wp_valid = BtbPlugin_logic_memWrite_valid;
  assign BtbPlugin_logic_memDp_wp_payload_address = BtbPlugin_logic_memWrite_payload_address;
  assign BtbPlugin_logic_memDp_wp_payload_data_0_hash = BtbPlugin_logic_memWrite_payload_data_0_hash;
  assign BtbPlugin_logic_memDp_wp_payload_data_0_sliceLow = BtbPlugin_logic_memWrite_payload_data_0_sliceLow;
  assign BtbPlugin_logic_memDp_wp_payload_data_0_pcTarget = BtbPlugin_logic_memWrite_payload_data_0_pcTarget;
  assign BtbPlugin_logic_memDp_wp_payload_data_0_isBranch = BtbPlugin_logic_memWrite_payload_data_0_isBranch;
  assign BtbPlugin_logic_memDp_wp_payload_data_0_isPush = BtbPlugin_logic_memWrite_payload_data_0_isPush;
  assign BtbPlugin_logic_memDp_wp_payload_data_0_isPop = BtbPlugin_logic_memWrite_payload_data_0_isPop;
  assign BtbPlugin_logic_memDp_wp_payload_mask = BtbPlugin_logic_memWrite_payload_mask;
  assign _zz_BtbPlugin_logic_memDp_rp_rsp_0_hash = BtbPlugin_logic_mem_spinal_port1[57 : 0];
  assign BtbPlugin_logic_memDp_rp_rsp_0_hash = _zz_BtbPlugin_logic_memDp_rp_rsp_0_hash[15 : 0];
  assign BtbPlugin_logic_memDp_rp_rsp_0_sliceLow = _zz_BtbPlugin_logic_memDp_rp_rsp_0_hash[16 : 16];
  assign BtbPlugin_logic_memDp_rp_rsp_0_pcTarget = _zz_BtbPlugin_logic_memDp_rp_rsp_0_hash[54 : 17];
  assign BtbPlugin_logic_memDp_rp_rsp_0_isBranch = _zz_BtbPlugin_logic_memDp_rp_rsp_0_hash[55];
  assign BtbPlugin_logic_memDp_rp_rsp_0_isPush = _zz_BtbPlugin_logic_memDp_rp_rsp_0_hash[56];
  assign BtbPlugin_logic_memDp_rp_rsp_0_isPop = _zz_BtbPlugin_logic_memDp_rp_rsp_0_hash[57];
  assign BtbPlugin_logic_memDp_rp_cmd_valid = BtbPlugin_logic_memRead_cmd_valid;
  assign BtbPlugin_logic_memDp_rp_cmd_payload = BtbPlugin_logic_memRead_cmd_payload;
  assign BtbPlugin_logic_memRead_rsp_0_hash = BtbPlugin_logic_memDp_rp_rsp_0_hash;
  assign BtbPlugin_logic_memRead_rsp_0_sliceLow = BtbPlugin_logic_memDp_rp_rsp_0_sliceLow;
  assign BtbPlugin_logic_memRead_rsp_0_pcTarget = BtbPlugin_logic_memDp_rp_rsp_0_pcTarget;
  assign BtbPlugin_logic_memRead_rsp_0_isBranch = BtbPlugin_logic_memDp_rp_rsp_0_isBranch;
  assign BtbPlugin_logic_memRead_rsp_0_isPush = BtbPlugin_logic_memDp_rp_rsp_0_isPush;
  assign BtbPlugin_logic_memRead_rsp_0_isPop = BtbPlugin_logic_memDp_rp_rsp_0_isPop;
  assign WhiteboxerPlugin_logic_fetch_fetchId = fetch_logic_ctrls_0_down_Fetch_ID;
  assign WhiteboxerPlugin_logic_decodes_0_fire = ((decode_ctrls_0_up_LANE_SEL_0 && decode_ctrls_0_up_isReady) && (! decode_ctrls_0_lane0_upIsCancel));
  assign when_CtrlLaneApi_l50 = (decode_ctrls_0_up_isReady || decode_ctrls_0_lane0_upIsCancel);
  assign WhiteboxerPlugin_logic_decodes_0_spawn = (decode_ctrls_0_up_LANE_SEL_0 && (! decode_ctrls_0_up_LANE_SEL_0_regNext));
  assign WhiteboxerPlugin_logic_decodes_0_pc = _zz_WhiteboxerPlugin_logic_decodes_0_pc;
  assign WhiteboxerPlugin_logic_decodes_0_fetchId = decode_ctrls_0_down_Fetch_ID_0;
  assign WhiteboxerPlugin_logic_decodes_0_decodeId = decode_ctrls_0_down_Decode_DOP_ID_0;
  always @(*) begin
    early0_EnvPlugin_logic_flushPort_valid = 1'b0;
    if(when_EnvPlugin_l119) begin
      early0_EnvPlugin_logic_flushPort_valid = 1'b1;
    end
  end

  assign early0_EnvPlugin_logic_flushPort_payload_uopId = execute_ctrl2_down_Decode_UOP_ID_lane0;
  assign early0_EnvPlugin_logic_flushPort_payload_self = 1'b0;
  always @(*) begin
    early0_EnvPlugin_logic_trapPort_valid = 1'b0;
    if(when_EnvPlugin_l119) begin
      early0_EnvPlugin_logic_trapPort_valid = 1'b1;
    end
  end

  always @(*) begin
    early0_EnvPlugin_logic_trapPort_payload_exception = 1'b1;
    case(execute_ctrl2_down_early0_EnvPlugin_OP_lane0)
      EnvPluginOp_EBREAK : begin
      end
      EnvPluginOp_ECALL : begin
      end
      EnvPluginOp_PRIV_RET : begin
        if(when_EnvPlugin_l86) begin
          early0_EnvPlugin_logic_trapPort_payload_exception = 1'b0;
        end
      end
      EnvPluginOp_WFI : begin
        if(when_EnvPlugin_l95) begin
          early0_EnvPlugin_logic_trapPort_payload_exception = 1'b0;
        end
      end
      EnvPluginOp_FENCE_I : begin
        early0_EnvPlugin_logic_trapPort_payload_exception = 1'b0;
      end
      default : begin
        if(when_EnvPlugin_l110) begin
          early0_EnvPlugin_logic_trapPort_payload_exception = 1'b0;
        end
      end
    endcase
  end

  assign MmuPlugin_logic_satpModeWrite = CsrAccessPlugin_bus_write_bits[63 : 60];
  assign FetchL1Plugin_pmaBuilder_addressBits = FetchL1Plugin_logic_ctrl_pmaPort_cmd_address;
  assign _zz_FetchL1Plugin_logic_ctrl_pmaPort_rsp_io = ((FetchL1Plugin_pmaBuilder_addressBits & 32'h0) == 32'h0);
  assign FetchL1Plugin_pmaBuilder_onTransfers_0_addressHit = _zz_FetchL1Plugin_pmaBuilder_onTransfers_0_addressHit[0];
  assign FetchL1Plugin_pmaBuilder_onTransfers_0_argsHit = (|1'b1);
  assign FetchL1Plugin_pmaBuilder_onTransfers_0_hit = (FetchL1Plugin_pmaBuilder_onTransfers_0_argsHit && FetchL1Plugin_pmaBuilder_onTransfers_0_addressHit);
  assign FetchL1Plugin_logic_ctrl_pmaPort_rsp_fault = (! ((|{((FetchL1Plugin_pmaBuilder_addressBits & 32'hf8000000) == 32'h80000000),((FetchL1Plugin_pmaBuilder_addressBits & 32'hf1000000) == 32'h0)}) && (|FetchL1Plugin_pmaBuilder_onTransfers_0_hit)));
  assign FetchL1Plugin_logic_ctrl_pmaPort_rsp_io = (! _zz_FetchL1Plugin_logic_ctrl_pmaPort_rsp_io_1[0]);
  assign FetchL1Axi4Plugin_logic_axi_ar_valid = FetchL1Plugin_logic_bus_cmd_valid;
  assign FetchL1Axi4Plugin_logic_axi_ar_payload_addr = FetchL1Plugin_logic_bus_cmd_payload_address;
  assign FetchL1Axi4Plugin_logic_axi_ar_payload_prot = 3'b110;
  assign FetchL1Axi4Plugin_logic_axi_ar_payload_cache = 4'b1111;
  assign FetchL1Axi4Plugin_logic_axi_ar_payload_len = 8'h07;
  assign FetchL1Axi4Plugin_logic_axi_ar_payload_size = 3'b011;
  assign FetchL1Axi4Plugin_logic_axi_ar_payload_burst = 2'b01;
  assign FetchL1Plugin_logic_bus_cmd_ready = FetchL1Axi4Plugin_logic_axi_ar_ready;
  assign FetchL1Plugin_logic_bus_rsp_valid = FetchL1Axi4Plugin_logic_axi_r_valid;
  assign FetchL1Plugin_logic_bus_rsp_payload_data = FetchL1Axi4Plugin_logic_axi_r_payload_data;
  assign FetchL1Plugin_logic_bus_rsp_payload_error = (! (FetchL1Axi4Plugin_logic_axi_r_payload_resp == 2'b00));
  assign FetchL1Axi4Plugin_logic_axi_r_ready = 1'b1;
  always @(*) begin
    DecoderPlugin_logic_forgetPort_valid = 1'b0;
    if(DecoderPlugin_logic_laneLogic_0_fixer_doIt) begin
      DecoderPlugin_logic_forgetPort_valid = 1'b1;
    end
  end

  always @(*) begin
    DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice = 39'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(DecoderPlugin_logic_laneLogic_0_fixer_doIt) begin
      DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice = (decode_ctrls_1_down_PC_0 + _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice);
    end
  end

  assign PerformanceCounterPlugin_logic_commitMask = PrivilegedPlugin_logic_harts_0_commitMask;
  assign when_PerformanceCounterPlugin_l45 = (|PerformanceCounterPlugin_logic_commitMask);
  assign PerformanceCounterPlugin_logic_commitCount = (_zz_PerformanceCounterPlugin_logic_commitCount - (PerformanceCounterPlugin_logic_ignoreNextCommit && (|PerformanceCounterPlugin_logic_commitMask)));
  assign PerformanceCounterPlugin_logic_counters_cycle_needFlush = PerformanceCounterPlugin_logic_counters_cycle_value[7];
  assign PerformanceCounterPlugin_logic_counters_instret_needFlush = PerformanceCounterPlugin_logic_counters_instret_value[7];
  assign PerformanceCounterPlugin_logic_eventCycles = 1'b1;
  assign PerformanceCounterPlugin_logic_eventInstructions_0 = _zz_PerformanceCounterPlugin_logic_eventInstructions_0[0];
  assign LsuPlugin_logic_cbmCsr_menvcfg_privLower = (PrivilegedPlugin_logic_harts_0_privilege < 2'b11);
  assign when_LsuPlugin_l226 = (LsuPlugin_logic_cbmCsr_menvcfg_privLower && (LsuPlugin_logic_cbmCsr_menvcfg_cbie == 2'b01));
  assign LsuPlugin_logic_cbmCsr_senvcfg_privLower = (PrivilegedPlugin_logic_harts_0_privilege < 2'b01);
  assign when_LsuPlugin_l226_1 = (LsuPlugin_logic_cbmCsr_senvcfg_privLower && (LsuPlugin_logic_cbmCsr_senvcfg_cbie == 2'b01));
  assign execute_ctrl0_down_AguPlugin_SIZE_lane0 = execute_ctrl0_down_Decode_UOP_lane0[13 : 12];
  assign LsuPlugin_logic_flusher_wantExit = 1'b0;
  always @(*) begin
    LsuPlugin_logic_flusher_wantStart = 1'b0;
    case(LsuPlugin_logic_flusher_stateReg)
      LsuPlugin_logic_flusher_CMD : begin
      end
      LsuPlugin_logic_flusher_COMPLETION : begin
      end
      default : begin
        LsuPlugin_logic_flusher_wantStart = 1'b1;
      end
    endcase
  end

  assign LsuPlugin_logic_flusher_wantKill = 1'b0;
  assign TrapPlugin_logic_lsuL1Invalidate_0_cmd_ready = LsuPlugin_logic_flusher_arbiter_io_inputs_0_ready;
  assign LsuPlugin_logic_flusher_inflight = (|{(execute_ctrl4_down_LsuL1_SEL_lane0 && execute_ctrl4_down_LsuL1_FLUSH_lane0),(execute_ctrl3_down_LsuL1_SEL_lane0 && execute_ctrl3_down_LsuL1_FLUSH_lane0)});
  always @(*) begin
    LsuPlugin_logic_flusher_arbiter_io_output_ready = 1'b0;
    case(LsuPlugin_logic_flusher_stateReg)
      LsuPlugin_logic_flusher_CMD : begin
      end
      LsuPlugin_logic_flusher_COMPLETION : begin
        if(when_LsuPlugin_l376) begin
          LsuPlugin_logic_flusher_arbiter_io_output_ready = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign PrivilegedPlugin_api_lsuTriggerBus_load = execute_ctrl3_down_LsuL1_LOAD_lane0;
  assign PrivilegedPlugin_api_lsuTriggerBus_store = execute_ctrl3_down_LsuL1_STORE_lane0;
  assign PrivilegedPlugin_api_lsuTriggerBus_virtual = execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0;
  assign PrivilegedPlugin_api_lsuTriggerBus_size = execute_ctrl3_down_LsuL1_SIZE_lane0;
  assign execute_ctrl3_down_LsuPlugin_logic_onTrigger_HIT_lane0 = 1'b0;
  assign execute_ctrl2_down_LsuPlugin_logic_FORCE_PHYSICAL_lane0 = (execute_ctrl2_down_LsuPlugin_logic_FROM_ACCESS_lane0 || execute_ctrl2_down_LsuPlugin_logic_FROM_WB_lane0);
  assign LsuPlugin_logic_onAddress0_ls_prefetchOp = execute_ctrl2_down_Decode_UOP_lane0[24 : 20];
  assign LsuPlugin_logic_onAddress0_ls_port_valid = (execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_down_AguPlugin_SEL_lane0);
  assign LsuPlugin_logic_onAddress0_ls_port_payload_address = _zz_LsuPlugin_logic_onAddress0_ls_port_payload_address[38:0];
  assign LsuPlugin_logic_onAddress0_ls_port_payload_size = execute_ctrl2_down_AguPlugin_SIZE_lane0;
  assign LsuPlugin_logic_onAddress0_ls_port_payload_load = execute_ctrl2_down_AguPlugin_LOAD_lane0;
  assign LsuPlugin_logic_onAddress0_ls_port_payload_store = execute_ctrl2_down_AguPlugin_STORE_lane0;
  assign LsuPlugin_logic_onAddress0_ls_port_payload_atomic = execute_ctrl2_down_AguPlugin_ATOMIC_lane0;
  assign LsuPlugin_logic_onAddress0_ls_port_payload_clean = (execute_ctrl2_down_AguPlugin_CLEAN_lane0 || (execute_ctrl2_down_AguPlugin_INVALIDATE_lane0 && LsuPlugin_logic_cbmCsr_invalIntoClean));
  assign LsuPlugin_logic_onAddress0_ls_port_payload_invalidate = execute_ctrl2_down_AguPlugin_INVALIDATE_lane0;
  assign LsuPlugin_logic_onAddress0_ls_port_payload_op = LsuL1CmdOpcode_LSU;
  assign LsuPlugin_logic_onAddress0_ls_port_fire = (LsuPlugin_logic_onAddress0_ls_port_valid && LsuPlugin_logic_onAddress0_ls_port_ready);
  assign LsuPlugin_logic_onAddress0_ls_port_payload_storeId = LsuPlugin_logic_onAddress0_ls_storeId;
  assign when_LsuPlugin_l264 = (|(LsuPlugin_logic_onAddress0_access_waiter_refill & (~ LsuL1_REFILL_BUSY)));
  assign LsuPlugin_logic_onAddress0_access_sbWaiter = 1'b0;
  assign _zz_MmuPlugin_logic_accessBus_cmd_ready = (! (LsuPlugin_logic_onAddress0_access_waiter_valid || LsuPlugin_logic_onAddress0_access_sbWaiter));
  assign MmuPlugin_logic_accessBus_cmd_haltWhen_valid = (MmuPlugin_logic_accessBus_cmd_valid && _zz_MmuPlugin_logic_accessBus_cmd_ready);
  assign MmuPlugin_logic_accessBus_cmd_ready = (MmuPlugin_logic_accessBus_cmd_haltWhen_ready && _zz_MmuPlugin_logic_accessBus_cmd_ready);
  assign MmuPlugin_logic_accessBus_cmd_haltWhen_payload_address = MmuPlugin_logic_accessBus_cmd_payload_address;
  assign MmuPlugin_logic_accessBus_cmd_haltWhen_payload_size = MmuPlugin_logic_accessBus_cmd_payload_size;
  assign LsuPlugin_logic_onAddress0_access_port_valid = MmuPlugin_logic_accessBus_cmd_haltWhen_valid;
  assign MmuPlugin_logic_accessBus_cmd_haltWhen_ready = LsuPlugin_logic_onAddress0_access_port_ready;
  assign LsuPlugin_logic_onAddress0_access_port_payload_address = {7'd0, MmuPlugin_logic_accessBus_cmd_payload_address};
  assign LsuPlugin_logic_onAddress0_access_port_payload_size = MmuPlugin_logic_accessBus_cmd_payload_size;
  assign LsuPlugin_logic_onAddress0_access_port_payload_load = 1'b1;
  assign LsuPlugin_logic_onAddress0_access_port_payload_store = 1'b0;
  assign LsuPlugin_logic_onAddress0_access_port_payload_atomic = 1'b0;
  assign LsuPlugin_logic_onAddress0_access_port_payload_clean = 1'b0;
  assign LsuPlugin_logic_onAddress0_access_port_payload_invalidate = 1'b0;
  assign LsuPlugin_logic_onAddress0_access_port_payload_op = LsuL1CmdOpcode_ACCESS_1;
  assign LsuPlugin_logic_onAddress0_access_port_payload_storeId = 12'h0;
  assign LsuPlugin_logic_onAddress0_flush_port_valid = ((LsuPlugin_logic_flusher_stateReg == LsuPlugin_logic_flusher_CMD) && (! LsuPlugin_logic_flusher_cmdCounter[6]));
  assign LsuPlugin_logic_onAddress0_flush_port_payload_address = {26'd0, _zz_LsuPlugin_logic_onAddress0_flush_port_payload_address};
  assign LsuPlugin_logic_onAddress0_flush_port_payload_size = 2'b00;
  assign LsuPlugin_logic_onAddress0_flush_port_payload_load = 1'b0;
  assign LsuPlugin_logic_onAddress0_flush_port_payload_store = 1'b0;
  assign LsuPlugin_logic_onAddress0_flush_port_payload_atomic = 1'b0;
  assign LsuPlugin_logic_onAddress0_flush_port_payload_clean = 1'b0;
  assign LsuPlugin_logic_onAddress0_flush_port_payload_invalidate = 1'b0;
  assign LsuPlugin_logic_onAddress0_flush_port_payload_op = LsuL1CmdOpcode_FLUSH;
  assign LsuPlugin_logic_onAddress0_flush_port_payload_storeId = 12'h0;
  assign LsuPlugin_logic_onAddress0_flush_port_fire = (LsuPlugin_logic_onAddress0_flush_port_valid && LsuPlugin_logic_onAddress0_flush_port_ready);
  assign LsuPlugin_logic_onAddress0_ls_port_ready = LsuPlugin_logic_onAddress0_arbiter_io_inputs_0_ready;
  assign LsuPlugin_logic_onAddress0_access_port_ready = LsuPlugin_logic_onAddress0_arbiter_io_inputs_1_ready;
  assign LsuPlugin_logic_onAddress0_flush_port_ready = LsuPlugin_logic_onAddress0_arbiter_io_inputs_2_ready;
  assign LsuPlugin_logic_onAddress0_arbiter_io_output_ready = (! execute_freeze_valid);
  assign execute_ctrl2_down_LsuL1_SEL_lane0 = LsuPlugin_logic_onAddress0_arbiter_io_output_valid;
  assign execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0 = LsuPlugin_logic_onAddress0_arbiter_io_output_payload_address;
  always @(*) begin
    _zz_execute_ctrl2_down_LsuL1_MASK_lane0 = 8'bxxxxxxxx;
    case(LsuPlugin_logic_onAddress0_arbiter_io_output_payload_size)
      2'b00 : begin
        _zz_execute_ctrl2_down_LsuL1_MASK_lane0 = 8'h01;
      end
      2'b01 : begin
        _zz_execute_ctrl2_down_LsuL1_MASK_lane0 = 8'h03;
      end
      2'b10 : begin
        _zz_execute_ctrl2_down_LsuL1_MASK_lane0 = 8'h0f;
      end
      default : begin
        _zz_execute_ctrl2_down_LsuL1_MASK_lane0 = 8'hff;
      end
    endcase
  end

  assign execute_ctrl2_down_LsuL1_MASK_lane0 = (_zz_execute_ctrl2_down_LsuL1_MASK_lane0 <<< LsuPlugin_logic_onAddress0_arbiter_io_output_payload_address[2 : 0]);
  assign execute_ctrl2_down_LsuL1_SIZE_lane0 = LsuPlugin_logic_onAddress0_arbiter_io_output_payload_size;
  assign execute_ctrl2_down_LsuL1_LOAD_lane0 = LsuPlugin_logic_onAddress0_arbiter_io_output_payload_load;
  assign execute_ctrl2_down_LsuL1_ATOMIC_lane0 = LsuPlugin_logic_onAddress0_arbiter_io_output_payload_atomic;
  assign execute_ctrl2_down_LsuL1_STORE_lane0 = LsuPlugin_logic_onAddress0_arbiter_io_output_payload_store;
  assign execute_ctrl2_down_LsuL1_CLEAN_lane0 = LsuPlugin_logic_onAddress0_arbiter_io_output_payload_clean;
  assign execute_ctrl2_down_LsuL1_INVALID_lane0 = LsuPlugin_logic_onAddress0_arbiter_io_output_payload_invalidate;
  assign execute_ctrl2_down_LsuL1_PREFETCH_lane0 = (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_op == LsuL1CmdOpcode_PREFETCH);
  assign execute_ctrl2_down_LsuL1_FLUSH_lane0 = (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_op == LsuL1CmdOpcode_FLUSH);
  assign execute_ctrl2_down_Decode_STORE_ID_lane0 = LsuPlugin_logic_onAddress0_arbiter_io_output_payload_storeId;
  assign execute_ctrl2_down_LsuPlugin_logic_FROM_ACCESS_lane0 = (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_op == LsuL1CmdOpcode_ACCESS_1);
  assign execute_ctrl2_down_LsuPlugin_logic_FROM_WB_lane0 = (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_op == LsuL1CmdOpcode_STORE_BUFFER);
  assign execute_ctrl2_down_LsuPlugin_logic_FROM_LSU_lane0 = (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_op == LsuL1CmdOpcode_LSU);
  assign execute_ctrl2_down_LsuPlugin_logic_FROM_PREFETCH_lane0 = (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_op == LsuL1CmdOpcode_PREFETCH);
  assign when_LsuPlugin_l529 = (! execute_ctrl2_down_LsuPlugin_logic_FROM_LSU_lane0);
  assign execute_ctrl3_down_LsuL1_PHYSICAL_ADDRESS_lane0 = execute_ctrl3_down_MMU_TRANSLATED_lane0;
  assign when_LsuPlugin_l557 = (execute_ctrl3_down_LsuPlugin_logic_FROM_LSU_lane0 && (! execute_ctrl3_up_LANE_SEL_lane0));
  assign when_LsuPlugin_l557_1 = (execute_ctrl4_down_LsuPlugin_logic_FROM_LSU_lane0 && (! execute_ctrl4_up_LANE_SEL_lane0));
  always @(*) begin
    execute_ctrl3_down_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0 = (|{((execute_ctrl3_down_LsuL1_SIZE_lane0 == 2'b11) && (execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[2 : 0] != 3'b000)),{((execute_ctrl3_down_LsuL1_SIZE_lane0 == 2'b10) && (execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[1 : 0] != 2'b00)),((execute_ctrl3_down_LsuL1_SIZE_lane0 == 2'b01) && (execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[0 : 0] != 1'b0))}});
    if(when_LsuPlugin_l565) begin
      execute_ctrl3_down_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0 = 1'b0;
    end
  end

  assign when_LsuPlugin_l565 = (execute_ctrl3_down_LsuL1_CLEAN_lane0 || execute_ctrl3_down_LsuL1_INVALID_lane0);
  assign execute_ctrl3_down_LsuPlugin_logic_preCtrl_IS_AMO_lane0 = (((execute_ctrl3_down_AguPlugin_SEL_lane0 && execute_ctrl3_down_LsuL1_ATOMIC_lane0) && execute_ctrl3_down_LsuL1_STORE_lane0) && execute_ctrl3_down_LsuL1_LOAD_lane0);
  assign LsuPlugin_logic_onPma_cached_cmd_address = execute_ctrl3_down_MMU_TRANSLATED_lane0;
  assign LsuPlugin_logic_onPma_cached_cmd_op[0] = execute_ctrl3_down_LsuL1_STORE_lane0;
  assign LsuPlugin_logic_onPma_io_cmd_address = execute_ctrl3_down_MMU_TRANSLATED_lane0;
  assign LsuPlugin_logic_onPma_io_cmd_size = execute_ctrl3_down_LsuL1_SIZE_lane0;
  assign LsuPlugin_logic_onPma_io_cmd_op[0] = execute_ctrl3_down_LsuL1_STORE_lane0;
  assign execute_ctrl3_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault = LsuPlugin_logic_onPma_cached_rsp_fault;
  assign execute_ctrl3_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_io = LsuPlugin_logic_onPma_cached_rsp_io;
  always @(*) begin
    execute_ctrl3_down_LsuPlugin_logic_onPma_IO_RSP_lane0_fault = LsuPlugin_logic_onPma_io_rsp_fault;
    if(when_LsuPlugin_l580) begin
      execute_ctrl3_down_LsuPlugin_logic_onPma_IO_RSP_lane0_fault = 1'b1;
    end
  end

  assign execute_ctrl3_down_LsuPlugin_logic_onPma_IO_RSP_lane0_io = LsuPlugin_logic_onPma_io_rsp_io;
  assign when_LsuPlugin_l580 = (execute_ctrl3_down_LsuL1_ATOMIC_lane0 || execute_ctrl3_down_LsuPlugin_logic_FROM_ACCESS_lane0);
  assign execute_ctrl3_down_LsuPlugin_logic_onPma_IO_lane0 = (((execute_ctrl3_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault && (! execute_ctrl3_down_LsuPlugin_logic_onPma_IO_RSP_lane0_fault)) && (! execute_ctrl3_down_LsuPlugin_logic_FENCE_lane0)) && (! execute_ctrl3_down_LsuPlugin_logic_FROM_PREFETCH_lane0));
  assign LsuPlugin_logic_onPma_addressExtension = (MmuPlugin_api_lsuTranslationEnable ? _zz_LsuPlugin_logic_onPma_addressExtension[38] : 1'b0);
  assign _zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0 = _zz__zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0;
  assign execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0 = (execute_ctrl3_down_LsuPlugin_logic_FROM_LSU_lane0 && (|{(_zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0[24] != LsuPlugin_logic_onPma_addressExtension),{(_zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0[23] != LsuPlugin_logic_onPma_addressExtension),{(_zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0[22] != LsuPlugin_logic_onPma_addressExtension),{(_zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0_1 != LsuPlugin_logic_onPma_addressExtension),{_zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0_2,{_zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0_3,_zz_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0_4}}}}}}));
  assign execute_ctrl3_down_LsuPlugin_logic_MMU_PAGE_FAULT_lane0 = (execute_ctrl3_down_MMU_PAGE_FAULT_lane0 || (execute_ctrl3_down_AguPlugin_STORE_lane0 ? (! execute_ctrl3_down_MMU_ALLOW_WRITE_lane0) : (! execute_ctrl3_down_MMU_ALLOW_READ_lane0)));
  assign execute_ctrl3_down_LsuPlugin_logic_MMU_FAILURE_lane0 = ((((execute_ctrl3_down_LsuPlugin_logic_MMU_PAGE_FAULT_lane0 || execute_ctrl3_down_MMU_ACCESS_FAULT_lane0) || execute_ctrl3_down_MMU_REFILL_lane0) || execute_ctrl3_down_MMU_HAZARD_lane0) || execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0);
  always @(*) begin
    LsuPlugin_logic_onCtrl_lsuTrap = 1'b0;
    if(LsuPlugin_logic_onCtrl_traps_accessFault) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b1;
    end
    if(LsuPlugin_logic_onCtrl_traps_l1Failed) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b1;
    end
    if(execute_ctrl4_down_LsuL1_CBM_REDO_lane0) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b1;
    end
    if(LsuPlugin_logic_onCtrl_traps_pmaFault) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b1;
    end
    if(execute_ctrl4_down_LsuPlugin_logic_MMU_PAGE_FAULT_lane0) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b1;
    end
    if(execute_ctrl4_down_MMU_ACCESS_FAULT_lane0) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b1;
    end
    if(execute_ctrl4_down_MMU_REFILL_lane0) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b1;
    end
    if(execute_ctrl4_down_MMU_HAZARD_lane0) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b1;
    end
    if(execute_ctrl4_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b1;
    end
    if(execute_ctrl4_down_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b1;
    end
    if(execute_ctrl4_down_LsuPlugin_logic_onTrigger_HIT_lane0) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b1;
    end
    if(when_LsuPlugin_l847) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b0;
    end
    if(when_LsuPlugin_l857) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b1;
    end
  end

  always @(*) begin
    LsuPlugin_logic_onCtrl_writeData = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    LsuPlugin_logic_onCtrl_writeData[63 : 0] = execute_ctrl4_up_integer_RS2_lane0;
    if(execute_ctrl4_down_LsuPlugin_logic_preCtrl_IS_AMO_lane0) begin
      LsuPlugin_logic_onCtrl_writeData[63 : 0] = LsuPlugin_logic_onCtrl_rva_aluBuffer;
    end
  end

  assign when_LsuPlugin_l608 = (((((! LsuPlugin_logic_onCtrl_lsuTrap) && (! execute_lane0_ctrls_4_upIsCancel)) && execute_ctrl4_down_LsuPlugin_logic_FROM_LSU_lane0) && (! execute_ctrl4_down_LsuL1_CLEAN_lane0)) && (! execute_ctrl4_down_LsuL1_INVALID_lane0));
  assign LsuPlugin_logic_onCtrl_io_doIt = ((execute_ctrl4_up_LANE_SEL_lane0 && execute_ctrl4_down_LsuL1_SEL_lane0) && execute_ctrl4_down_LsuPlugin_logic_onPma_IO_lane0);
  assign LsuPlugin_logic_bus_cmd_fire = (LsuPlugin_logic_bus_cmd_valid && LsuPlugin_logic_bus_cmd_ready);
  assign when_LsuPlugin_l612 = (! execute_freeze_valid);
  assign LsuPlugin_logic_bus_cmd_valid = (((LsuPlugin_logic_onCtrl_io_doItReg && (! LsuPlugin_logic_onCtrl_io_cmdSent)) && LsuPlugin_logic_onCtrl_io_allowIt) && (! LsuPlugin_logic_onCtrl_io_tooEarly));
  assign LsuPlugin_logic_bus_cmd_payload_write = execute_ctrl4_down_LsuL1_STORE_lane0;
  assign LsuPlugin_logic_bus_cmd_payload_address = execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0;
  assign LsuPlugin_logic_bus_cmd_payload_data = execute_ctrl4_down_LsuL1_WRITE_DATA_lane0;
  assign LsuPlugin_logic_bus_cmd_payload_size = execute_ctrl4_down_LsuL1_SIZE_lane0;
  assign LsuPlugin_logic_bus_cmd_payload_mask = execute_ctrl4_down_LsuL1_MASK_lane0;
  assign LsuPlugin_logic_bus_cmd_payload_io = 1'b1;
  assign LsuPlugin_logic_bus_cmd_payload_fromHart = 1'b1;
  assign LsuPlugin_logic_bus_cmd_payload_uopId = execute_ctrl4_down_Decode_UOP_ID_lane0;
  assign LsuPlugin_logic_bus_rsp_toStream_valid = LsuPlugin_logic_bus_rsp_valid;
  assign LsuPlugin_logic_bus_rsp_toStream_payload_error = LsuPlugin_logic_bus_rsp_payload_error;
  assign LsuPlugin_logic_bus_rsp_toStream_payload_data = LsuPlugin_logic_bus_rsp_payload_data;
  assign LsuPlugin_logic_onCtrl_io_rsp_fire = (LsuPlugin_logic_onCtrl_io_rsp_valid && LsuPlugin_logic_onCtrl_io_rsp_ready);
  assign LsuPlugin_logic_bus_rsp_toStream_ready = (! LsuPlugin_logic_bus_rsp_toStream_rValid);
  assign LsuPlugin_logic_onCtrl_io_rsp_valid = LsuPlugin_logic_bus_rsp_toStream_rValid;
  assign LsuPlugin_logic_onCtrl_io_rsp_payload_error = LsuPlugin_logic_bus_rsp_toStream_rData_error;
  assign LsuPlugin_logic_onCtrl_io_rsp_payload_data = LsuPlugin_logic_bus_rsp_toStream_rData_data;
  assign LsuPlugin_logic_onCtrl_io_rsp_ready = (! execute_freeze_valid);
  assign LsuPlugin_logic_onCtrl_io_freezeIt = (LsuPlugin_logic_onCtrl_io_doIt && (LsuPlugin_logic_onCtrl_io_tooEarly || ((! LsuPlugin_logic_onCtrl_io_rsp_valid) && LsuPlugin_logic_onCtrl_io_allowIt)));
  assign LsuPlugin_logic_onCtrl_loadData_input = (LsuPlugin_logic_onCtrl_io_cmdSent ? LsuPlugin_logic_onCtrl_io_rsp_payload_data : execute_ctrl4_down_LsuL1_READ_DATA_lane0);
  assign LsuPlugin_logic_onCtrl_loadData_splitted_0 = LsuPlugin_logic_onCtrl_loadData_input[7 : 0];
  assign LsuPlugin_logic_onCtrl_loadData_splitted_1 = LsuPlugin_logic_onCtrl_loadData_input[15 : 8];
  assign LsuPlugin_logic_onCtrl_loadData_splitted_2 = LsuPlugin_logic_onCtrl_loadData_input[23 : 16];
  assign LsuPlugin_logic_onCtrl_loadData_splitted_3 = LsuPlugin_logic_onCtrl_loadData_input[31 : 24];
  assign LsuPlugin_logic_onCtrl_loadData_splitted_4 = LsuPlugin_logic_onCtrl_loadData_input[39 : 32];
  assign LsuPlugin_logic_onCtrl_loadData_splitted_5 = LsuPlugin_logic_onCtrl_loadData_input[47 : 40];
  assign LsuPlugin_logic_onCtrl_loadData_splitted_6 = LsuPlugin_logic_onCtrl_loadData_input[55 : 48];
  assign LsuPlugin_logic_onCtrl_loadData_splitted_7 = LsuPlugin_logic_onCtrl_loadData_input[63 : 56];
  always @(*) begin
    LsuPlugin_logic_onCtrl_loadData_shifted[7 : 0] = _zz_LsuPlugin_logic_onCtrl_loadData_shifted;
    LsuPlugin_logic_onCtrl_loadData_shifted[15 : 8] = _zz_LsuPlugin_logic_onCtrl_loadData_shifted_2;
    LsuPlugin_logic_onCtrl_loadData_shifted[23 : 16] = _zz_LsuPlugin_logic_onCtrl_loadData_shifted_4;
    LsuPlugin_logic_onCtrl_loadData_shifted[31 : 24] = _zz_LsuPlugin_logic_onCtrl_loadData_shifted_6;
    LsuPlugin_logic_onCtrl_loadData_shifted[39 : 32] = LsuPlugin_logic_onCtrl_loadData_splitted_4;
    LsuPlugin_logic_onCtrl_loadData_shifted[47 : 40] = LsuPlugin_logic_onCtrl_loadData_splitted_5;
    LsuPlugin_logic_onCtrl_loadData_shifted[55 : 48] = LsuPlugin_logic_onCtrl_loadData_splitted_6;
    LsuPlugin_logic_onCtrl_loadData_shifted[63 : 56] = LsuPlugin_logic_onCtrl_loadData_splitted_7;
  end

  assign execute_ctrl4_down_LsuPlugin_logic_onCtrl_loadData_RESULT_lane0 = LsuPlugin_logic_onCtrl_loadData_shifted;
  assign LsuPlugin_logic_onCtrl_storeData_mapping_0_1 = {8{LsuPlugin_logic_onCtrl_writeData[7 : 0]}};
  assign LsuPlugin_logic_onCtrl_storeData_mapping_1_1 = {4{LsuPlugin_logic_onCtrl_writeData[15 : 0]}};
  assign LsuPlugin_logic_onCtrl_storeData_mapping_2_1 = {2{LsuPlugin_logic_onCtrl_writeData[31 : 0]}};
  assign LsuPlugin_logic_onCtrl_storeData_mapping_3_1 = {1{LsuPlugin_logic_onCtrl_writeData[63 : 0]}};
  always @(*) begin
    _zz_execute_ctrl4_down_LsuL1_WRITE_DATA_lane0 = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(execute_ctrl4_down_LsuL1_SIZE_lane0)
      2'b00 : begin
        _zz_execute_ctrl4_down_LsuL1_WRITE_DATA_lane0 = LsuPlugin_logic_onCtrl_storeData_mapping_0_1;
      end
      2'b01 : begin
        _zz_execute_ctrl4_down_LsuL1_WRITE_DATA_lane0 = LsuPlugin_logic_onCtrl_storeData_mapping_1_1;
      end
      2'b10 : begin
        _zz_execute_ctrl4_down_LsuL1_WRITE_DATA_lane0 = LsuPlugin_logic_onCtrl_storeData_mapping_2_1;
      end
      default : begin
        _zz_execute_ctrl4_down_LsuL1_WRITE_DATA_lane0 = LsuPlugin_logic_onCtrl_storeData_mapping_3_1;
      end
    endcase
  end

  assign execute_ctrl4_down_LsuL1_WRITE_DATA_lane0 = _zz_execute_ctrl4_down_LsuL1_WRITE_DATA_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_onCtrl_SC_MISS_lane0 = LsuPlugin_logic_onCtrl_scMiss;
  assign _zz_LsuPlugin_logic_onCtrl_rva_alu_compare = execute_ctrl4_down_Decode_UOP_lane0[31 : 29];
  assign _zz_LsuPlugin_logic_onCtrl_rva_alu_selectRf = execute_ctrl4_down_Decode_UOP_lane0[27];
  assign when_Rvi_l230 = (execute_ctrl4_down_LsuL1_SIZE_lane0 == 2'b10);
  assign LsuPlugin_logic_onCtrl_rva_alu_compare = _zz_LsuPlugin_logic_onCtrl_rva_alu_compare[2];
  assign LsuPlugin_logic_onCtrl_rva_alu_unsigned = _zz_LsuPlugin_logic_onCtrl_rva_alu_compare[1];
  assign LsuPlugin_logic_onCtrl_rva_alu_addSub = _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub;
  always @(*) begin
    LsuPlugin_logic_onCtrl_rva_alu_less = ((execute_ctrl4_up_integer_RS2_lane0[63] == LsuPlugin_logic_onCtrl_rva_srcBuffer[63]) ? LsuPlugin_logic_onCtrl_rva_alu_addSub[63] : (LsuPlugin_logic_onCtrl_rva_alu_unsigned ? LsuPlugin_logic_onCtrl_rva_srcBuffer[63] : execute_ctrl4_up_integer_RS2_lane0[63]));
    if(when_Rvi_l230) begin
      LsuPlugin_logic_onCtrl_rva_alu_less = ((execute_ctrl4_up_integer_RS2_lane0[31] == LsuPlugin_logic_onCtrl_rva_srcBuffer[31]) ? LsuPlugin_logic_onCtrl_rva_alu_addSub[31] : (LsuPlugin_logic_onCtrl_rva_alu_unsigned ? LsuPlugin_logic_onCtrl_rva_srcBuffer[31] : execute_ctrl4_up_integer_RS2_lane0[31]));
    end
  end

  assign LsuPlugin_logic_onCtrl_rva_alu_selectRf = (_zz_LsuPlugin_logic_onCtrl_rva_alu_selectRf ? 1'b1 : (_zz_LsuPlugin_logic_onCtrl_rva_alu_compare[0] ^ LsuPlugin_logic_onCtrl_rva_alu_less));
  assign switch_Misc_l245 = (_zz_LsuPlugin_logic_onCtrl_rva_alu_compare | {_zz_LsuPlugin_logic_onCtrl_rva_alu_selectRf,2'b00});
  always @(*) begin
    case(switch_Misc_l245)
      3'b000 : begin
        LsuPlugin_logic_onCtrl_rva_alu_raw = LsuPlugin_logic_onCtrl_rva_alu_addSub;
      end
      3'b001 : begin
        LsuPlugin_logic_onCtrl_rva_alu_raw = (execute_ctrl4_up_integer_RS2_lane0 ^ LsuPlugin_logic_onCtrl_rva_srcBuffer);
      end
      3'b010 : begin
        LsuPlugin_logic_onCtrl_rva_alu_raw = (execute_ctrl4_up_integer_RS2_lane0 | LsuPlugin_logic_onCtrl_rva_srcBuffer);
      end
      3'b011 : begin
        LsuPlugin_logic_onCtrl_rva_alu_raw = (execute_ctrl4_up_integer_RS2_lane0 & LsuPlugin_logic_onCtrl_rva_srcBuffer);
      end
      default : begin
        LsuPlugin_logic_onCtrl_rva_alu_raw = (LsuPlugin_logic_onCtrl_rva_alu_selectRf ? execute_ctrl4_up_integer_RS2_lane0 : LsuPlugin_logic_onCtrl_rva_srcBuffer);
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_onCtrl_rva_alu_result = LsuPlugin_logic_onCtrl_rva_alu_raw;
    if(when_Rvi_l230) begin
      LsuPlugin_logic_onCtrl_rva_alu_result[63 : 32] = (LsuPlugin_logic_onCtrl_rva_alu_raw[31] ? 32'hffffffff : 32'h0);
    end
  end

  assign LsuPlugin_logic_onCtrl_rva_delay_0 = _zz_LsuPlugin_logic_onCtrl_rva_delay_0;
  assign LsuPlugin_logic_onCtrl_rva_delay_1 = _zz_LsuPlugin_logic_onCtrl_rva_delay_1;
  assign LsuPlugin_logic_onCtrl_rva_freezeIt = ((execute_ctrl4_up_LANE_SEL_lane0 && execute_ctrl4_down_LsuPlugin_logic_preCtrl_IS_AMO_lane0) && (|{LsuPlugin_logic_onCtrl_rva_delay_1,LsuPlugin_logic_onCtrl_rva_delay_0}));
  always @(*) begin
    LsuPlugin_logic_onCtrl_rva_lrsc_capture = 1'b0;
    if(when_LsuPlugin_l697) begin
      if(!execute_ctrl4_down_LsuL1_STORE_lane0) begin
        if(execute_ctrl4_down_LsuL1_ATOMIC_lane0) begin
          LsuPlugin_logic_onCtrl_rva_lrsc_capture = 1'b1;
        end
      end
    end
  end

  assign when_LsuPlugin_l697 = ((((((! execute_freeze_valid) && execute_ctrl4_up_LANE_SEL_lane0) && execute_ctrl4_down_LsuPlugin_logic_FROM_LSU_lane0) && execute_ctrl4_down_LsuL1_SEL_lane0) && (! LsuPlugin_logic_onCtrl_lsuTrap)) && (! execute_ctrl4_down_LsuPlugin_logic_onPma_IO_lane0));
  assign LsuPlugin_logic_onCtrl_scMiss = (! LsuPlugin_logic_onCtrl_rva_lrsc_reserved);
  assign LsuL1_lockPort_valid = LsuPlugin_logic_onCtrl_rva_lrsc_reserved;
  assign LsuL1_lockPort_address = LsuPlugin_logic_onCtrl_rva_lrsc_address;
  assign when_LsuPlugin_l709 = ((! LsuPlugin_logic_onCtrl_rva_lrsc_age[5]) && (! execute_freeze_valid));
  assign when_LsuPlugin_l716 = ((LsuPlugin_logic_onCtrl_rva_lrsc_age[5] || LsuPlugin_logic_onCtrl_io_cmdSent) || LsuL1Plugin_logic_slotsFreezeHazard);
  assign when_LsuPlugin_l720 = (LsuPlugin_logic_onCtrl_rva_lrsc_capture && (LsuPlugin_logic_onCtrl_rva_lrsc_reserved || (6'h08 <= LsuPlugin_logic_onCtrl_rva_lrsc_age)));
  always @(*) begin
    LsuPlugin_logic_flushPort_valid = 1'b0;
    if(when_LsuPlugin_l908) begin
      if(LsuPlugin_logic_onCtrl_lsuTrap) begin
        LsuPlugin_logic_flushPort_valid = 1'b1;
      end
    end
  end

  assign LsuPlugin_logic_flushPort_payload_uopId = execute_ctrl4_down_Decode_UOP_ID_lane0;
  assign LsuPlugin_logic_flushPort_payload_self = 1'b0;
  always @(*) begin
    LsuPlugin_logic_trapPort_valid = 1'b0;
    if(when_LsuPlugin_l908) begin
      if(LsuPlugin_logic_onCtrl_lsuTrap) begin
        LsuPlugin_logic_trapPort_valid = 1'b1;
      end
    end
  end

  assign LsuPlugin_logic_trapPort_payload_tval = execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0;
  always @(*) begin
    LsuPlugin_logic_trapPort_payload_exception = 1'bx;
    if(LsuPlugin_logic_onCtrl_traps_accessFault) begin
      LsuPlugin_logic_trapPort_payload_exception = 1'b1;
    end
    if(LsuPlugin_logic_onCtrl_traps_l1Failed) begin
      LsuPlugin_logic_trapPort_payload_exception = 1'b0;
    end
    if(execute_ctrl4_down_LsuL1_CBM_REDO_lane0) begin
      LsuPlugin_logic_trapPort_payload_exception = 1'b0;
    end
    if(LsuPlugin_logic_onCtrl_traps_pmaFault) begin
      LsuPlugin_logic_trapPort_payload_exception = 1'b1;
    end
    if(execute_ctrl4_down_LsuPlugin_logic_MMU_PAGE_FAULT_lane0) begin
      LsuPlugin_logic_trapPort_payload_exception = 1'b1;
    end
    if(execute_ctrl4_down_MMU_ACCESS_FAULT_lane0) begin
      LsuPlugin_logic_trapPort_payload_exception = 1'b1;
    end
    if(execute_ctrl4_down_MMU_REFILL_lane0) begin
      LsuPlugin_logic_trapPort_payload_exception = 1'b0;
    end
    if(execute_ctrl4_down_MMU_HAZARD_lane0) begin
      LsuPlugin_logic_trapPort_payload_exception = 1'b0;
    end
    if(execute_ctrl4_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0) begin
      LsuPlugin_logic_trapPort_payload_exception = 1'b1;
    end
    if(execute_ctrl4_down_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0) begin
      LsuPlugin_logic_trapPort_payload_exception = 1'b1;
    end
    if(execute_ctrl4_down_LsuPlugin_logic_onTrigger_HIT_lane0) begin
      LsuPlugin_logic_trapPort_payload_exception = 1'b0;
    end
    if(when_LsuPlugin_l857) begin
      LsuPlugin_logic_trapPort_payload_exception = 1'b0;
    end
  end

  always @(*) begin
    LsuPlugin_logic_trapPort_payload_code = 4'bxxxx;
    if(LsuPlugin_logic_onCtrl_traps_accessFault) begin
      LsuPlugin_logic_trapPort_payload_code = 4'b0101;
      if(execute_ctrl4_down_LsuL1_STORE_lane0) begin
        LsuPlugin_logic_trapPort_payload_code[1] = 1'b1;
      end
    end
    if(LsuPlugin_logic_onCtrl_traps_l1Failed) begin
      LsuPlugin_logic_trapPort_payload_code = 4'b0100;
    end
    if(execute_ctrl4_down_LsuL1_CBM_REDO_lane0) begin
      LsuPlugin_logic_trapPort_payload_code = 4'b0100;
    end
    if(LsuPlugin_logic_onCtrl_traps_pmaFault) begin
      LsuPlugin_logic_trapPort_payload_code = 4'b0101;
      if(execute_ctrl4_down_LsuL1_STORE_lane0) begin
        LsuPlugin_logic_trapPort_payload_code[1] = 1'b1;
      end
    end
    if(execute_ctrl4_down_LsuPlugin_logic_MMU_PAGE_FAULT_lane0) begin
      LsuPlugin_logic_trapPort_payload_code = 4'b1101;
      if(execute_ctrl4_down_LsuL1_STORE_lane0) begin
        LsuPlugin_logic_trapPort_payload_code[1] = 1'b1;
      end
    end
    if(execute_ctrl4_down_MMU_ACCESS_FAULT_lane0) begin
      LsuPlugin_logic_trapPort_payload_code = 4'b0101;
      if(execute_ctrl4_down_LsuL1_STORE_lane0) begin
        LsuPlugin_logic_trapPort_payload_code[1] = 1'b1;
      end
    end
    if(execute_ctrl4_down_MMU_REFILL_lane0) begin
      LsuPlugin_logic_trapPort_payload_code = 4'b0111;
    end
    if(execute_ctrl4_down_MMU_HAZARD_lane0) begin
      LsuPlugin_logic_trapPort_payload_code = 4'b0100;
    end
    if(execute_ctrl4_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0) begin
      LsuPlugin_logic_trapPort_payload_code = 4'b0101;
      if(execute_ctrl4_down_AguPlugin_STORE_lane0) begin
        LsuPlugin_logic_trapPort_payload_code[1] = 1'b1;
      end
      if(when_LsuPlugin_l820) begin
        LsuPlugin_logic_trapPort_payload_code[3] = 1'b1;
      end
    end
    if(execute_ctrl4_down_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0) begin
      LsuPlugin_logic_trapPort_payload_code = {1'd0, _zz_LsuPlugin_logic_trapPort_payload_code};
    end
    if(execute_ctrl4_down_LsuPlugin_logic_onTrigger_HIT_lane0) begin
      LsuPlugin_logic_trapPort_payload_code = 4'b0011;
    end
    if(when_LsuPlugin_l857) begin
      LsuPlugin_logic_trapPort_payload_code = 4'b0100;
    end
  end

  always @(*) begin
    LsuPlugin_logic_trapPort_payload_arg = 3'b000;
    LsuPlugin_logic_trapPort_payload_arg[1 : 0] = (execute_ctrl4_down_LsuL1_STORE_lane0 ? 2'b01 : 2'b00);
    LsuPlugin_logic_trapPort_payload_arg[2 : 2] = 1'b1;
  end

  assign LsuPlugin_logic_onCtrl_traps_accessFault = ((execute_ctrl4_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault ? (LsuPlugin_logic_onCtrl_io_rsp_valid && LsuPlugin_logic_onCtrl_io_rsp_payload_error) : execute_ctrl4_down_LsuL1_FAULT_lane0) || execute_ctrl4_down_LsuPlugin_logic_pmpPort_ACCESS_FAULT_lane0);
  assign LsuPlugin_logic_onCtrl_traps_l1Failed = (execute_ctrl4_down_LsuL1_SEL_lane0 && ((! execute_ctrl4_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault) && (execute_ctrl4_down_LsuL1_HAZARD_lane0 || ((execute_ctrl4_down_LsuL1_MISS_lane0 || execute_ctrl4_down_LsuL1_MISS_UNIQUE_lane0) && (execute_ctrl4_down_LsuL1_LOAD_lane0 || execute_ctrl4_down_LsuL1_STORE_lane0)))));
  assign LsuPlugin_logic_onCtrl_traps_pmaFault = (execute_ctrl4_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault && execute_ctrl4_down_LsuPlugin_logic_onPma_IO_RSP_lane0_fault);
  assign when_LsuPlugin_l820 = (! execute_ctrl4_down_MMU_BYPASS_TRANSLATION_lane0);
  assign when_LsuPlugin_l847 = (execute_ctrl4_down_LsuPlugin_logic_FENCE_lane0 || execute_ctrl4_down_LsuPlugin_logic_FROM_PREFETCH_lane0);
  assign LsuPlugin_logic_onCtrl_fenceTrap_enable = 1'b0;
  always @(*) begin
    LsuPlugin_logic_onCtrl_fenceTrap_doIt = ((execute_ctrl4_down_LsuL1_ATOMIC_lane0 || execute_ctrl4_down_LsuPlugin_logic_FENCE_lane0) && LsuPlugin_logic_onCtrl_fenceTrap_enable);
    if(LsuPlugin_logic_onCtrl_cmbTrap_valid) begin
      LsuPlugin_logic_onCtrl_fenceTrap_doIt = 1'b1;
    end
  end

  assign when_LsuPlugin_l855 = (! execute_freeze_valid);
  assign when_LsuPlugin_l857 = (LsuPlugin_logic_onCtrl_fenceTrap_doIt || LsuPlugin_logic_onCtrl_fenceTrap_doItReg);
  assign when_LsuPlugin_l897 = (! execute_freeze_valid);
  assign LsuPlugin_logic_onCtrl_cmbTrap_pending = (LsuPlugin_logic_onCtrl_cmbTrap_cmbTrigger || (|LsuPlugin_logic_onCtrl_cmbTrap_pendingWritebacks));
  assign LsuPlugin_logic_onCtrl_cmbTrap_valid = (((execute_ctrl4_down_LsuL1_ATOMIC_lane0 || execute_ctrl4_down_LsuPlugin_logic_FENCE_lane0) || execute_ctrl4_down_LsuL1_LOAD_lane0) && LsuPlugin_logic_onCtrl_cmbTrap_pending);
  assign when_LsuPlugin_l908 = (execute_ctrl4_up_LANE_SEL_lane0 && execute_ctrl4_down_AguPlugin_SEL_lane0);
  assign LsuPlugin_logic_onCtrl_mmuNeeded = (execute_ctrl4_down_LsuPlugin_logic_FROM_LSU_lane0 || execute_ctrl4_down_LsuPlugin_logic_FROM_PREFETCH_lane0);
  assign execute_ctrl4_down_LsuL1_ABORD_lane0 = (|{(execute_ctrl4_down_LsuPlugin_logic_FROM_LSU_lane0 && (LsuPlugin_logic_onCtrl_fenceTrap_doIt || LsuPlugin_logic_onCtrl_fenceTrap_doItReg)),{(LsuPlugin_logic_onCtrl_mmuNeeded && execute_ctrl4_down_LsuPlugin_logic_MMU_FAILURE_lane0),{(execute_ctrl4_down_LsuPlugin_logic_FROM_LSU_lane0 && ((_zz_execute_ctrl4_down_LsuL1_ABORD_lane0 || execute_lane0_ctrls_4_upIsCancel) || execute_ctrl4_down_LsuPlugin_logic_FENCE_lane0)),{((! execute_ctrl4_down_LsuL1_FLUSH_lane0) && execute_ctrl4_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault),{execute_ctrl4_down_LsuL1_FLUSH_HAZARD_lane0,execute_ctrl4_down_LsuL1_HAZARD_lane0}}}}});
  assign execute_ctrl4_down_LsuL1_SKIP_WRITE_lane0 = (|{((execute_ctrl4_down_LsuL1_ATOMIC_lane0 && (! execute_ctrl4_down_LsuL1_LOAD_lane0)) && LsuPlugin_logic_onCtrl_scMiss),{execute_ctrl4_down_LsuPlugin_logic_FROM_PREFETCH_lane0,{(execute_ctrl4_down_LsuPlugin_logic_FROM_LSU_lane0 && (execute_ctrl4_down_LsuPlugin_logic_onTrigger_HIT_lane0 || execute_ctrl4_down_LsuPlugin_logic_pmpPort_ACCESS_FAULT_lane0)),{execute_ctrl4_down_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0,{execute_ctrl4_down_LsuL1_FAULT_lane0,(execute_ctrl4_down_LsuL1_MISS_lane0 || execute_ctrl4_down_LsuL1_MISS_UNIQUE_lane0)}}}}});
  assign when_LsuPlugin_l949 = ((execute_ctrl4_down_LsuL1_SEL_lane0 && execute_ctrl4_down_LsuL1_FLUSH_lane0) && ((execute_ctrl4_down_LsuL1_FLUSH_HIT_lane0 || execute_ctrl4_down_LsuL1_HAZARD_lane0) || execute_ctrl4_down_LsuL1_FLUSH_HAZARD_lane0));
  assign MmuPlugin_logic_accessBus_rsp_valid = ((execute_ctrl4_down_LsuL1_SEL_lane0 && execute_ctrl4_down_LsuPlugin_logic_FROM_ACCESS_lane0) && (! execute_freeze_valid));
  assign MmuPlugin_logic_accessBus_rsp_payload_data = execute_ctrl4_down_LsuPlugin_logic_onCtrl_loadData_RESULT_lane0;
  always @(*) begin
    MmuPlugin_logic_accessBus_rsp_payload_error = (execute_ctrl4_down_LsuL1_FAULT_lane0 || execute_ctrl4_down_LsuPlugin_logic_pmpPort_ACCESS_FAULT_lane0);
    if(LsuPlugin_logic_onCtrl_traps_pmaFault) begin
      MmuPlugin_logic_accessBus_rsp_payload_error = 1'b1;
    end
  end

  always @(*) begin
    MmuPlugin_logic_accessBus_rsp_payload_redo = LsuPlugin_logic_onCtrl_traps_l1Failed;
    if(LsuPlugin_logic_onCtrl_traps_pmaFault) begin
      MmuPlugin_logic_accessBus_rsp_payload_redo = 1'b0;
    end
  end

  assign MmuPlugin_logic_accessBus_rsp_payload_waitAny = 1'b0;
  assign when_LsuPlugin_l986 = (MmuPlugin_logic_accessBus_rsp_valid && MmuPlugin_logic_accessBus_rsp_payload_redo);
  assign when_LsuPlugin_l268 = (|execute_ctrl4_down_LsuL1_WAIT_REFILL_lane0);
  assign when_LsuPlugin_l264_1 = (|(LsuPlugin_logic_onCtrl_hartRegulation_refill & (~ LsuL1_REFILL_BUSY)));
  assign when_LsuPlugin_l993 = ((((((execute_ctrl4_up_LANE_SEL_lane0 && execute_ctrl4_down_AguPlugin_SEL_lane0) && (! execute_ctrl4_down_LsuPlugin_logic_FROM_PREFETCH_lane0)) && (! execute_ctrl4_down_LsuPlugin_logic_onPma_IO_lane0)) && (! execute_ctrl4_down_LsuPlugin_logic_FENCE_lane0)) && 1'b1) && ((execute_ctrl4_down_LsuL1_HAZARD_lane0 || execute_ctrl4_down_LsuL1_MISS_lane0) || execute_ctrl4_down_LsuL1_MISS_UNIQUE_lane0));
  assign when_LsuPlugin_l268_1 = (|execute_ctrl4_down_LsuL1_WAIT_REFILL_lane0);
  assign LsuPlugin_logic_onCtrl_commitProbeReq = ((((((((((execute_ctrl4_down_LANE_SEL_lane0 && execute_ctrl4_down_isReady) && (! execute_lane0_ctrls_4_downIsCancel)) && execute_ctrl4_down_AguPlugin_SEL_lane0) && execute_ctrl4_down_LsuPlugin_logic_FROM_LSU_lane0) && (execute_ctrl4_down_LsuL1_LOAD_lane0 || execute_ctrl4_down_LsuL1_STORE_lane0)) && (! execute_ctrl4_down_LsuL1_PREFETCH_lane0)) && (! execute_ctrl4_down_LsuL1_ATOMIC_lane0)) && (! execute_ctrl4_down_LsuL1_FLUSH_lane0)) && (! execute_ctrl4_down_LsuL1_CLEAN_lane0)) && (! execute_ctrl4_down_LsuL1_INVALID_lane0));
  assign LsuPlugin_logic_commitProbe_valid = (LsuPlugin_logic_onCtrl_commitProbeReq && (! LsuPlugin_logic_onCtrl_commitProbeToken));
  assign LsuPlugin_logic_commitProbe_payload_address = execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0;
  assign LsuPlugin_logic_commitProbe_payload_load = execute_ctrl4_down_LsuL1_LOAD_lane0;
  assign LsuPlugin_logic_commitProbe_payload_store = execute_ctrl4_down_LsuL1_STORE_lane0;
  assign LsuPlugin_logic_commitProbe_payload_trap = LsuPlugin_logic_onCtrl_lsuTrap;
  assign LsuPlugin_logic_commitProbe_payload_miss = ((((execute_ctrl4_down_LsuL1_MISS_lane0 || execute_ctrl4_down_LsuL1_MISS_UNIQUE_lane0) || execute_ctrl4_down_LsuL1_HAZARD_lane0) && (! execute_ctrl4_down_LsuPlugin_logic_MMU_FAILURE_lane0)) && 1'b1);
  assign LsuPlugin_logic_commitProbe_payload_io = execute_ctrl4_down_LsuPlugin_logic_onPma_IO_lane0;
  assign LsuPlugin_logic_commitProbe_payload_prefetchFailed = execute_ctrl4_down_LsuPlugin_logic_FROM_PREFETCH_lane0;
  assign LsuPlugin_logic_commitProbe_payload_pc = execute_ctrl4_down_PC_lane0;
  assign LsuPlugin_logic_iwb_valid = (execute_ctrl4_down_AguPlugin_SEL_lane0 && (! execute_ctrl4_down_AguPlugin_FLOAT_lane0));
  always @(*) begin
    LsuPlugin_logic_iwb_payload = execute_ctrl4_down_LsuPlugin_logic_onCtrl_loadData_RESULT_lane0;
    if(when_LsuPlugin_l1018) begin
      LsuPlugin_logic_iwb_payload[0] = execute_ctrl4_down_LsuPlugin_logic_onCtrl_SC_MISS_lane0;
      LsuPlugin_logic_iwb_payload[7 : 1] = 7'h0;
    end
  end

  assign when_LsuPlugin_l1018 = (execute_ctrl4_down_LsuL1_ATOMIC_lane0 && (! execute_ctrl4_down_LsuL1_LOAD_lane0));
  assign LsuPlugin_logic_onWb_storeFire = ((((((execute_ctrl4_down_LANE_SEL_lane0 && execute_ctrl4_down_isReady) && (! execute_lane0_ctrls_4_downIsCancel)) && execute_ctrl4_down_AguPlugin_SEL_lane0) && execute_ctrl4_down_LsuL1_STORE_lane0) && (! execute_ctrl4_down_LsuPlugin_logic_onPma_IO_lane0)) && (! execute_ctrl4_down_LsuPlugin_logic_FROM_PREFETCH_lane0));
  assign LsuPlugin_logic_onWb_storeBroadcast = (((((((execute_ctrl4_down_isReady && execute_ctrl4_down_LsuL1_SEL_lane0) && execute_ctrl4_down_LsuL1_STORE_lane0) && (! execute_ctrl4_down_LsuL1_ABORD_lane0)) && (! execute_ctrl4_down_LsuL1_SKIP_WRITE_lane0)) && (! execute_ctrl4_down_LsuL1_MISS_lane0)) && (! execute_ctrl4_down_LsuL1_MISS_UNIQUE_lane0)) && (! execute_ctrl4_down_LsuL1_HAZARD_lane0));
  always @(*) begin
    _zz_execute_ctrl1_down_early0_SrcPlugin_SRC1_lane0 = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(execute_ctrl1_down_early0_SrcPlugin_logic_SRC1_CTRL_lane0)
      1'b0 : begin
        _zz_execute_ctrl1_down_early0_SrcPlugin_SRC1_lane0 = execute_ctrl1_down_integer_RS1_lane0;
      end
      default : begin
        _zz_execute_ctrl1_down_early0_SrcPlugin_SRC1_lane0 = {{32{_zz__zz_execute_ctrl1_down_early0_SrcPlugin_SRC1_lane0[31]}}, _zz__zz_execute_ctrl1_down_early0_SrcPlugin_SRC1_lane0};
      end
    endcase
  end

  assign execute_ctrl1_down_early0_SrcPlugin_SRC1_lane0 = _zz_execute_ctrl1_down_early0_SrcPlugin_SRC1_lane0;
  always @(*) begin
    _zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0 = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(execute_ctrl1_down_early0_SrcPlugin_logic_SRC2_CTRL_lane0)
      2'b00 : begin
        _zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0 = execute_ctrl1_down_integer_RS2_lane0;
      end
      2'b01 : begin
        _zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0 = {{52{_zz__zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0[11]}}, _zz__zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0};
      end
      2'b10 : begin
        _zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0 = {{25{_zz__zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0_1[38]}}, _zz__zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0_1};
      end
      default : begin
        _zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0 = {{52{_zz__zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0_2[11]}}, _zz__zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0_2};
      end
    endcase
  end

  assign execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0 = _zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0;
  always @(*) begin
    early0_SrcPlugin_logic_addsub_combined_rs2Patched = execute_ctrl2_down_early0_SrcPlugin_SRC2_lane0;
    if(execute_ctrl2_down_SrcStageables_REVERT_lane0) begin
      early0_SrcPlugin_logic_addsub_combined_rs2Patched = (~ execute_ctrl2_down_early0_SrcPlugin_SRC2_lane0);
    end
    if(execute_ctrl2_down_SrcStageables_ZERO_lane0) begin
      early0_SrcPlugin_logic_addsub_combined_rs2Patched = 64'h0;
    end
  end

  assign execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0 = ($signed(_zz_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0) + $signed(_zz_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0_1));
  assign execute_ctrl2_down_early0_SrcPlugin_LESS_lane0 = ((execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[63] == execute_ctrl2_down_early0_SrcPlugin_SRC2_lane0[63]) ? execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0[63] : (execute_ctrl2_down_SrcStageables_UNSIGNED_lane0 ? execute_ctrl2_down_early0_SrcPlugin_SRC2_lane0[63] : execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[63]));
  assign lane0_IntFormatPlugin_logic_stages_0_hits = {early0_BarrelShifterPlugin_logic_wb_valid,early0_IntAluPlugin_logic_wb_valid};
  assign lane0_IntFormatPlugin_logic_stages_0_wb_valid = (execute_ctrl2_up_LANE_SEL_lane0 && (|lane0_IntFormatPlugin_logic_stages_0_hits));
  assign lane0_IntFormatPlugin_logic_stages_0_raw = ((lane0_IntFormatPlugin_logic_stages_0_hits[0] ? early0_IntAluPlugin_logic_wb_payload : 64'h0) | (lane0_IntFormatPlugin_logic_stages_0_hits[1] ? early0_BarrelShifterPlugin_logic_wb_payload : 64'h0));
  always @(*) begin
    lane0_IntFormatPlugin_logic_stages_0_wb_payload = lane0_IntFormatPlugin_logic_stages_0_raw;
    if(lane0_IntFormatPlugin_logic_stages_0_segments_0_doIt) begin
      lane0_IntFormatPlugin_logic_stages_0_wb_payload[63 : 32] = {32{lane0_IntFormatPlugin_logic_stages_0_segments_0_sign_value}};
    end
  end

  assign lane0_IntFormatPlugin_logic_stages_0_segments_0_sign_sels_0 = lane0_IntFormatPlugin_logic_stages_0_raw[31];
  always @(*) begin
    _zz_lane0_IntFormatPlugin_logic_stages_0_segments_0_sign_value = 1'bx;
    case(execute_ctrl2_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0)
      2'b10 : begin
        _zz_lane0_IntFormatPlugin_logic_stages_0_segments_0_sign_value = lane0_IntFormatPlugin_logic_stages_0_segments_0_sign_sels_0;
      end
      default : begin
      end
    endcase
  end

  assign lane0_IntFormatPlugin_logic_stages_0_segments_0_sign_value = (execute_ctrl2_down_lane0_IntFormatPlugin_logic_SIGNED_lane0 && _zz_lane0_IntFormatPlugin_logic_stages_0_segments_0_sign_value);
  assign lane0_IntFormatPlugin_logic_stages_0_segments_0_doIt = (execute_ctrl2_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0 < 2'b11);
  assign lane0_IntFormatPlugin_logic_stages_1_hits = {LsuPlugin_logic_iwb_valid,early0_MulPlugin_logic_formatBus_valid};
  assign lane0_IntFormatPlugin_logic_stages_1_wb_valid = (execute_ctrl4_up_LANE_SEL_lane0 && (|lane0_IntFormatPlugin_logic_stages_1_hits));
  assign lane0_IntFormatPlugin_logic_stages_1_raw = ((lane0_IntFormatPlugin_logic_stages_1_hits[0] ? early0_MulPlugin_logic_formatBus_payload : 64'h0) | (lane0_IntFormatPlugin_logic_stages_1_hits[1] ? LsuPlugin_logic_iwb_payload : 64'h0));
  always @(*) begin
    lane0_IntFormatPlugin_logic_stages_1_wb_payload = lane0_IntFormatPlugin_logic_stages_1_raw;
    if(lane0_IntFormatPlugin_logic_stages_1_segments_0_doIt) begin
      lane0_IntFormatPlugin_logic_stages_1_wb_payload[15 : 8] = {8{lane0_IntFormatPlugin_logic_stages_1_segments_0_sign_value}};
    end
    if(lane0_IntFormatPlugin_logic_stages_1_segments_1_doIt) begin
      lane0_IntFormatPlugin_logic_stages_1_wb_payload[31 : 16] = {16{lane0_IntFormatPlugin_logic_stages_1_segments_1_sign_value}};
    end
    if(lane0_IntFormatPlugin_logic_stages_1_segments_2_doIt) begin
      lane0_IntFormatPlugin_logic_stages_1_wb_payload[63 : 32] = {32{lane0_IntFormatPlugin_logic_stages_1_segments_2_sign_value}};
    end
  end

  assign lane0_IntFormatPlugin_logic_stages_1_segments_0_sign_sels_0 = lane0_IntFormatPlugin_logic_stages_1_raw[7];
  always @(*) begin
    _zz_lane0_IntFormatPlugin_logic_stages_1_segments_0_sign_value = 1'bx;
    case(execute_ctrl4_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0)
      2'b00 : begin
        _zz_lane0_IntFormatPlugin_logic_stages_1_segments_0_sign_value = lane0_IntFormatPlugin_logic_stages_1_segments_0_sign_sels_0;
      end
      default : begin
      end
    endcase
  end

  assign lane0_IntFormatPlugin_logic_stages_1_segments_0_sign_value = (execute_ctrl4_down_lane0_IntFormatPlugin_logic_SIGNED_lane0 && _zz_lane0_IntFormatPlugin_logic_stages_1_segments_0_sign_value);
  assign lane0_IntFormatPlugin_logic_stages_1_segments_0_doIt = (execute_ctrl4_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0 < 2'b01);
  assign lane0_IntFormatPlugin_logic_stages_1_segments_1_sign_sels_0 = lane0_IntFormatPlugin_logic_stages_1_raw[7];
  assign lane0_IntFormatPlugin_logic_stages_1_segments_1_sign_sels_1 = lane0_IntFormatPlugin_logic_stages_1_raw[15];
  always @(*) begin
    _zz_lane0_IntFormatPlugin_logic_stages_1_segments_1_sign_value = 1'bx;
    case(execute_ctrl4_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0)
      2'b00 : begin
        _zz_lane0_IntFormatPlugin_logic_stages_1_segments_1_sign_value = lane0_IntFormatPlugin_logic_stages_1_segments_1_sign_sels_0;
      end
      2'b01 : begin
        _zz_lane0_IntFormatPlugin_logic_stages_1_segments_1_sign_value = lane0_IntFormatPlugin_logic_stages_1_segments_1_sign_sels_1;
      end
      default : begin
      end
    endcase
  end

  assign lane0_IntFormatPlugin_logic_stages_1_segments_1_sign_value = (execute_ctrl4_down_lane0_IntFormatPlugin_logic_SIGNED_lane0 && _zz_lane0_IntFormatPlugin_logic_stages_1_segments_1_sign_value);
  assign lane0_IntFormatPlugin_logic_stages_1_segments_1_doIt = (execute_ctrl4_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0 < 2'b10);
  assign lane0_IntFormatPlugin_logic_stages_1_segments_2_sign_sels_0 = lane0_IntFormatPlugin_logic_stages_1_raw[31];
  assign lane0_IntFormatPlugin_logic_stages_1_segments_2_sign_sels_1 = lane0_IntFormatPlugin_logic_stages_1_raw[7];
  assign lane0_IntFormatPlugin_logic_stages_1_segments_2_sign_sels_2 = lane0_IntFormatPlugin_logic_stages_1_raw[15];
  always @(*) begin
    _zz_lane0_IntFormatPlugin_logic_stages_1_segments_2_sign_value = 1'bx;
    case(execute_ctrl4_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0)
      2'b10 : begin
        _zz_lane0_IntFormatPlugin_logic_stages_1_segments_2_sign_value = lane0_IntFormatPlugin_logic_stages_1_segments_2_sign_sels_0;
      end
      2'b00 : begin
        _zz_lane0_IntFormatPlugin_logic_stages_1_segments_2_sign_value = lane0_IntFormatPlugin_logic_stages_1_segments_2_sign_sels_1;
      end
      2'b01 : begin
        _zz_lane0_IntFormatPlugin_logic_stages_1_segments_2_sign_value = lane0_IntFormatPlugin_logic_stages_1_segments_2_sign_sels_2;
      end
      default : begin
      end
    endcase
  end

  assign lane0_IntFormatPlugin_logic_stages_1_segments_2_sign_value = (execute_ctrl4_down_lane0_IntFormatPlugin_logic_SIGNED_lane0 && _zz_lane0_IntFormatPlugin_logic_stages_1_segments_2_sign_value);
  assign lane0_IntFormatPlugin_logic_stages_1_segments_2_doIt = (execute_ctrl4_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0 < 2'b11);
  assign lane0_IntFormatPlugin_logic_stages_2_hits = {CsrAccessPlugin_logic_wbWi_valid,early0_DivPlugin_logic_formatBus_valid};
  assign lane0_IntFormatPlugin_logic_stages_2_wb_valid = (execute_ctrl3_up_LANE_SEL_lane0 && (|lane0_IntFormatPlugin_logic_stages_2_hits));
  assign lane0_IntFormatPlugin_logic_stages_2_raw = ((lane0_IntFormatPlugin_logic_stages_2_hits[0] ? early0_DivPlugin_logic_formatBus_payload : 64'h0) | (lane0_IntFormatPlugin_logic_stages_2_hits[1] ? CsrAccessPlugin_logic_wbWi_payload : 64'h0));
  always @(*) begin
    lane0_IntFormatPlugin_logic_stages_2_wb_payload = lane0_IntFormatPlugin_logic_stages_2_raw;
    if(lane0_IntFormatPlugin_logic_stages_2_segments_0_doIt) begin
      lane0_IntFormatPlugin_logic_stages_2_wb_payload[63 : 32] = {32{lane0_IntFormatPlugin_logic_stages_2_segments_0_sign_value}};
    end
  end

  assign lane0_IntFormatPlugin_logic_stages_2_segments_0_sign_sels_0 = lane0_IntFormatPlugin_logic_stages_2_raw[31];
  always @(*) begin
    _zz_lane0_IntFormatPlugin_logic_stages_2_segments_0_sign_value = 1'bx;
    case(execute_ctrl3_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0)
      2'b10 : begin
        _zz_lane0_IntFormatPlugin_logic_stages_2_segments_0_sign_value = lane0_IntFormatPlugin_logic_stages_2_segments_0_sign_sels_0;
      end
      default : begin
      end
    endcase
  end

  assign lane0_IntFormatPlugin_logic_stages_2_segments_0_sign_value = (execute_ctrl3_down_lane0_IntFormatPlugin_logic_SIGNED_lane0 && _zz_lane0_IntFormatPlugin_logic_stages_2_segments_0_sign_value);
  assign lane0_IntFormatPlugin_logic_stages_2_segments_0_doIt = (execute_ctrl3_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0 < 2'b11);
  always @(*) begin
    case(execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0)
      BranchPlugin_BranchCtrlEnum_JALR : begin
        early0_BranchPlugin_pcCalc_target_a = execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[38:0];
      end
      default : begin
        early0_BranchPlugin_pcCalc_target_a = execute_ctrl2_down_PC_lane0;
      end
    endcase
  end

  always @(*) begin
    case(execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0)
      BranchPlugin_BranchCtrlEnum_JAL : begin
        early0_BranchPlugin_pcCalc_target_b = {{43{_zz_early0_BranchPlugin_pcCalc_target_b[20]}}, _zz_early0_BranchPlugin_pcCalc_target_b};
      end
      BranchPlugin_BranchCtrlEnum_JALR : begin
        early0_BranchPlugin_pcCalc_target_b = {{52{_zz_early0_BranchPlugin_pcCalc_target_b_1[11]}}, _zz_early0_BranchPlugin_pcCalc_target_b_1};
      end
      default : begin
        early0_BranchPlugin_pcCalc_target_b = {{51{_zz_early0_BranchPlugin_pcCalc_target_b_2[12]}}, _zz_early0_BranchPlugin_pcCalc_target_b_2};
      end
    endcase
  end

  assign early0_BranchPlugin_pcCalc_slices = ({1'b0,execute_ctrl2_down_Decode_INSTRUCTION_SLICE_COUNT_lane0} + {1'b0,1'b1});
  always @(*) begin
    execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0 = _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0[38:0];
    execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0[0] = 1'b0;
  end

  assign execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0 = (execute_ctrl2_down_PC_lane0 + _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0);
  assign execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0 = (execute_ctrl2_down_PC_lane0 + _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0);
  assign AlignerPlugin_logic_maskGen_frontMasks_0 = 2'b11;
  assign AlignerPlugin_logic_maskGen_frontMasks_1 = 2'b10;
  assign AlignerPlugin_logic_maskGen_backMasks_0 = 2'b01;
  assign AlignerPlugin_logic_maskGen_backMasks_1 = 2'b11;
  assign fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK = (_zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK & ((! fetch_logic_ctrls_2_down_Prediction_WORD_JUMPED) ? 2'b11 : _zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK_2));
  assign fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_LAST = ((fetch_logic_ctrls_2_up_isValid && fetch_logic_ctrls_2_down_Prediction_WORD_JUMPED) ? _zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_LAST : 2'b00);
  assign AlignerPlugin_logic_slicesInstructions_0 = {AlignerPlugin_logic_slices_data_1,AlignerPlugin_logic_slices_data_0};
  assign AlignerPlugin_logic_slicesInstructions_1 = {AlignerPlugin_logic_slices_data_2,AlignerPlugin_logic_slices_data_1};
  assign AlignerPlugin_logic_slicesInstructions_2 = {AlignerPlugin_logic_slices_data_3,AlignerPlugin_logic_slices_data_2};
  assign AlignerPlugin_logic_slicesInstructions_3 = {16'd0, AlignerPlugin_logic_slices_data_3};
  always @(*) begin
    AlignerPlugin_logic_scanners_0_usageMask = 4'b0000;
    AlignerPlugin_logic_scanners_0_usageMask[0] = AlignerPlugin_logic_scanners_0_checker_0_required;
    AlignerPlugin_logic_scanners_0_usageMask[1] = AlignerPlugin_logic_scanners_0_checker_1_required;
  end

  assign AlignerPlugin_logic_scanners_0_checker_0_required = 1'b1;
  assign AlignerPlugin_logic_scanners_0_checker_0_last = (AlignerPlugin_logic_slices_data_0[1 : 0] != 2'b11);
  assign AlignerPlugin_logic_scanners_0_checker_0_redo = ((AlignerPlugin_logic_scanners_0_checker_0_required && AlignerPlugin_logic_slices_last[0]) && (! AlignerPlugin_logic_scanners_0_checker_0_last));
  assign AlignerPlugin_logic_scanners_0_checker_0_present = AlignerPlugin_logic_slices_mask[0];
  assign AlignerPlugin_logic_scanners_0_checker_0_valid = AlignerPlugin_logic_scanners_0_checker_0_present;
  assign AlignerPlugin_logic_scanners_0_checker_1_required = (AlignerPlugin_logic_slices_data_0[1 : 0] == 2'b11);
  assign AlignerPlugin_logic_scanners_0_checker_1_last = (AlignerPlugin_logic_slices_data_0[1 : 0] == 2'b11);
  assign AlignerPlugin_logic_scanners_0_checker_1_redo = ((AlignerPlugin_logic_scanners_0_checker_1_required && AlignerPlugin_logic_slices_last[1]) && (! AlignerPlugin_logic_scanners_0_checker_1_last));
  assign AlignerPlugin_logic_scanners_0_checker_1_present = AlignerPlugin_logic_slices_mask[1];
  assign AlignerPlugin_logic_scanners_0_checker_1_valid = (AlignerPlugin_logic_scanners_0_checker_1_present || (! AlignerPlugin_logic_scanners_0_checker_1_required));
  assign AlignerPlugin_logic_scanners_0_redo = (|{AlignerPlugin_logic_scanners_0_checker_1_redo,AlignerPlugin_logic_scanners_0_checker_0_redo});
  assign AlignerPlugin_logic_scanners_0_valid = (AlignerPlugin_logic_scanners_0_checker_0_valid && ((&AlignerPlugin_logic_scanners_0_checker_1_valid) || (|{AlignerPlugin_logic_scanners_0_checker_1_redo,AlignerPlugin_logic_scanners_0_checker_0_redo})));
  always @(*) begin
    AlignerPlugin_logic_scanners_1_usageMask = 4'b0000;
    AlignerPlugin_logic_scanners_1_usageMask[1] = AlignerPlugin_logic_scanners_1_checker_0_required;
    AlignerPlugin_logic_scanners_1_usageMask[2] = AlignerPlugin_logic_scanners_1_checker_1_required;
  end

  assign AlignerPlugin_logic_scanners_1_checker_0_required = 1'b1;
  assign AlignerPlugin_logic_scanners_1_checker_0_last = (AlignerPlugin_logic_slices_data_1[1 : 0] != 2'b11);
  assign AlignerPlugin_logic_scanners_1_checker_0_redo = ((AlignerPlugin_logic_scanners_1_checker_0_required && AlignerPlugin_logic_slices_last[1]) && (! AlignerPlugin_logic_scanners_1_checker_0_last));
  assign AlignerPlugin_logic_scanners_1_checker_0_present = AlignerPlugin_logic_slices_mask[1];
  assign AlignerPlugin_logic_scanners_1_checker_0_valid = AlignerPlugin_logic_scanners_1_checker_0_present;
  assign AlignerPlugin_logic_scanners_1_checker_1_required = (AlignerPlugin_logic_slices_data_1[1 : 0] == 2'b11);
  assign AlignerPlugin_logic_scanners_1_checker_1_last = (AlignerPlugin_logic_slices_data_1[1 : 0] == 2'b11);
  assign AlignerPlugin_logic_scanners_1_checker_1_redo = ((AlignerPlugin_logic_scanners_1_checker_1_required && AlignerPlugin_logic_slices_last[2]) && (! AlignerPlugin_logic_scanners_1_checker_1_last));
  assign AlignerPlugin_logic_scanners_1_checker_1_present = AlignerPlugin_logic_slices_mask[2];
  assign AlignerPlugin_logic_scanners_1_checker_1_valid = (AlignerPlugin_logic_scanners_1_checker_1_present || (! AlignerPlugin_logic_scanners_1_checker_1_required));
  assign AlignerPlugin_logic_scanners_1_redo = (|{AlignerPlugin_logic_scanners_1_checker_1_redo,AlignerPlugin_logic_scanners_1_checker_0_redo});
  assign AlignerPlugin_logic_scanners_1_valid = (AlignerPlugin_logic_scanners_1_checker_0_valid && ((&AlignerPlugin_logic_scanners_1_checker_1_valid) || (|{AlignerPlugin_logic_scanners_1_checker_1_redo,AlignerPlugin_logic_scanners_1_checker_0_redo})));
  always @(*) begin
    AlignerPlugin_logic_scanners_2_usageMask = 4'b0000;
    AlignerPlugin_logic_scanners_2_usageMask[2] = AlignerPlugin_logic_scanners_2_checker_0_required;
    AlignerPlugin_logic_scanners_2_usageMask[3] = AlignerPlugin_logic_scanners_2_checker_1_required;
  end

  assign AlignerPlugin_logic_scanners_2_checker_0_required = 1'b1;
  assign AlignerPlugin_logic_scanners_2_checker_0_last = (AlignerPlugin_logic_slices_data_2[1 : 0] != 2'b11);
  assign AlignerPlugin_logic_scanners_2_checker_0_redo = ((AlignerPlugin_logic_scanners_2_checker_0_required && AlignerPlugin_logic_slices_last[2]) && (! AlignerPlugin_logic_scanners_2_checker_0_last));
  assign AlignerPlugin_logic_scanners_2_checker_0_present = AlignerPlugin_logic_slices_mask[2];
  assign AlignerPlugin_logic_scanners_2_checker_0_valid = AlignerPlugin_logic_scanners_2_checker_0_present;
  assign AlignerPlugin_logic_scanners_2_checker_1_required = (AlignerPlugin_logic_slices_data_2[1 : 0] == 2'b11);
  assign AlignerPlugin_logic_scanners_2_checker_1_last = (AlignerPlugin_logic_slices_data_2[1 : 0] == 2'b11);
  assign AlignerPlugin_logic_scanners_2_checker_1_redo = ((AlignerPlugin_logic_scanners_2_checker_1_required && AlignerPlugin_logic_slices_last[3]) && (! AlignerPlugin_logic_scanners_2_checker_1_last));
  assign AlignerPlugin_logic_scanners_2_checker_1_present = AlignerPlugin_logic_slices_mask[3];
  assign AlignerPlugin_logic_scanners_2_checker_1_valid = (AlignerPlugin_logic_scanners_2_checker_1_present || (! AlignerPlugin_logic_scanners_2_checker_1_required));
  assign AlignerPlugin_logic_scanners_2_redo = (|{AlignerPlugin_logic_scanners_2_checker_1_redo,AlignerPlugin_logic_scanners_2_checker_0_redo});
  assign AlignerPlugin_logic_scanners_2_valid = (AlignerPlugin_logic_scanners_2_checker_0_valid && ((&AlignerPlugin_logic_scanners_2_checker_1_valid) || (|{AlignerPlugin_logic_scanners_2_checker_1_redo,AlignerPlugin_logic_scanners_2_checker_0_redo})));
  always @(*) begin
    AlignerPlugin_logic_scanners_3_usageMask = 4'b0000;
    AlignerPlugin_logic_scanners_3_usageMask[3] = AlignerPlugin_logic_scanners_3_checker_0_required;
  end

  assign AlignerPlugin_logic_scanners_3_checker_0_required = 1'b1;
  assign AlignerPlugin_logic_scanners_3_checker_0_last = (AlignerPlugin_logic_slices_data_3[1 : 0] != 2'b11);
  assign AlignerPlugin_logic_scanners_3_checker_0_redo = ((AlignerPlugin_logic_scanners_3_checker_0_required && AlignerPlugin_logic_slices_last[3]) && (! AlignerPlugin_logic_scanners_3_checker_0_last));
  assign AlignerPlugin_logic_scanners_3_checker_0_present = AlignerPlugin_logic_slices_mask[3];
  assign AlignerPlugin_logic_scanners_3_checker_0_valid = AlignerPlugin_logic_scanners_3_checker_0_present;
  assign AlignerPlugin_logic_scanners_3_checker_1_required = (AlignerPlugin_logic_slices_data_3[1 : 0] == 2'b11);
  assign AlignerPlugin_logic_scanners_3_checker_1_last = (AlignerPlugin_logic_slices_data_3[1 : 0] == 2'b11);
  assign AlignerPlugin_logic_scanners_3_checker_1_redo = 1'b0;
  assign AlignerPlugin_logic_scanners_3_checker_1_present = 1'b0;
  assign AlignerPlugin_logic_scanners_3_checker_1_valid = (AlignerPlugin_logic_scanners_3_checker_1_present || (! AlignerPlugin_logic_scanners_3_checker_1_required));
  assign AlignerPlugin_logic_scanners_3_redo = (|{AlignerPlugin_logic_scanners_3_checker_1_redo,AlignerPlugin_logic_scanners_3_checker_0_redo});
  assign AlignerPlugin_logic_scanners_3_valid = (AlignerPlugin_logic_scanners_3_checker_0_valid && ((&AlignerPlugin_logic_scanners_3_checker_1_valid) || (|{AlignerPlugin_logic_scanners_3_checker_1_redo,AlignerPlugin_logic_scanners_3_checker_0_redo})));
  assign AlignerPlugin_logic_usedMask_0 = 4'b0000;
  assign AlignerPlugin_logic_extractors_0_first = 1'b1;
  assign AlignerPlugin_logic_extractors_0_usableMask = {(AlignerPlugin_logic_scanners_3_valid && (! AlignerPlugin_logic_usedMask_0[3])),{(AlignerPlugin_logic_scanners_2_valid && (! AlignerPlugin_logic_usedMask_0[2])),{(AlignerPlugin_logic_scanners_1_valid && (! AlignerPlugin_logic_usedMask_0[1])),(AlignerPlugin_logic_scanners_0_valid && (! AlignerPlugin_logic_usedMask_0[0]))}}};
  assign _zz_AlignerPlugin_logic_extractors_0_usableMask_bools_0 = AlignerPlugin_logic_extractors_0_usableMask;
  assign AlignerPlugin_logic_extractors_0_usableMask_bools_0 = _zz_AlignerPlugin_logic_extractors_0_usableMask_bools_0[0];
  assign AlignerPlugin_logic_extractors_0_usableMask_bools_1 = _zz_AlignerPlugin_logic_extractors_0_usableMask_bools_0[1];
  assign AlignerPlugin_logic_extractors_0_usableMask_bools_2 = _zz_AlignerPlugin_logic_extractors_0_usableMask_bools_0[2];
  assign AlignerPlugin_logic_extractors_0_usableMask_bools_3 = _zz_AlignerPlugin_logic_extractors_0_usableMask_bools_0[3];
  always @(*) begin
    _zz_AlignerPlugin_logic_extractors_0_slicesOh[0] = (AlignerPlugin_logic_extractors_0_usableMask_bools_0 && (! 1'b0));
    _zz_AlignerPlugin_logic_extractors_0_slicesOh[1] = (AlignerPlugin_logic_extractors_0_usableMask_bools_1 && (! AlignerPlugin_logic_extractors_0_usableMask_bools_0));
    _zz_AlignerPlugin_logic_extractors_0_slicesOh[2] = (AlignerPlugin_logic_extractors_0_usableMask_bools_2 && (! AlignerPlugin_logic_extractors_0_usableMask_range_0_to_1));
    _zz_AlignerPlugin_logic_extractors_0_slicesOh[3] = (AlignerPlugin_logic_extractors_0_usableMask_bools_3 && (! AlignerPlugin_logic_extractors_0_usableMask_range_0_to_2));
  end

  assign AlignerPlugin_logic_extractors_0_usableMask_range_0_to_1 = (|{AlignerPlugin_logic_extractors_0_usableMask_bools_1,AlignerPlugin_logic_extractors_0_usableMask_bools_0});
  assign AlignerPlugin_logic_extractors_0_usableMask_range_0_to_2 = (|{AlignerPlugin_logic_extractors_0_usableMask_bools_2,{AlignerPlugin_logic_extractors_0_usableMask_bools_1,AlignerPlugin_logic_extractors_0_usableMask_bools_0}});
  assign AlignerPlugin_logic_extractors_0_slicesOh = _zz_AlignerPlugin_logic_extractors_0_slicesOh;
  assign _zz_AlignerPlugin_logic_extractors_0_redo = AlignerPlugin_logic_extractors_0_slicesOh[0];
  assign _zz_AlignerPlugin_logic_extractors_0_redo_1 = AlignerPlugin_logic_extractors_0_slicesOh[1];
  assign _zz_AlignerPlugin_logic_extractors_0_redo_2 = AlignerPlugin_logic_extractors_0_slicesOh[2];
  assign _zz_AlignerPlugin_logic_extractors_0_redo_3 = AlignerPlugin_logic_extractors_0_slicesOh[3];
  always @(*) begin
    AlignerPlugin_logic_extractors_0_redo = _zz_AlignerPlugin_logic_extractors_0_redo_4[0];
    if(when_AlignerPlugin_l160) begin
      AlignerPlugin_logic_extractors_0_redo = 1'b0;
    end
  end

  assign AlignerPlugin_logic_extractors_0_localMask = (((_zz_AlignerPlugin_logic_extractors_0_redo ? {AlignerPlugin_logic_scanners_0_checker_1_required,AlignerPlugin_logic_scanners_0_checker_0_required} : 2'b00) | (_zz_AlignerPlugin_logic_extractors_0_redo_1 ? {AlignerPlugin_logic_scanners_1_checker_1_required,AlignerPlugin_logic_scanners_1_checker_0_required} : 2'b00)) | ((_zz_AlignerPlugin_logic_extractors_0_redo_2 ? {AlignerPlugin_logic_scanners_2_checker_1_required,AlignerPlugin_logic_scanners_2_checker_0_required} : 2'b00) | (_zz_AlignerPlugin_logic_extractors_0_redo_3 ? {AlignerPlugin_logic_scanners_3_checker_1_required,AlignerPlugin_logic_scanners_3_checker_0_required} : 2'b00)));
  assign AlignerPlugin_logic_extractors_0_usageMask = (((_zz_AlignerPlugin_logic_extractors_0_redo ? AlignerPlugin_logic_scanners_0_usageMask : 4'b0000) | (_zz_AlignerPlugin_logic_extractors_0_redo_1 ? AlignerPlugin_logic_scanners_1_usageMask : 4'b0000)) | ((_zz_AlignerPlugin_logic_extractors_0_redo_2 ? AlignerPlugin_logic_scanners_2_usageMask : 4'b0000) | (_zz_AlignerPlugin_logic_extractors_0_redo_3 ? AlignerPlugin_logic_scanners_3_usageMask : 4'b0000)));
  assign AlignerPlugin_logic_usedMask_1 = (AlignerPlugin_logic_usedMask_0 | AlignerPlugin_logic_extractors_0_usageMask);
  always @(*) begin
    AlignerPlugin_logic_extractors_0_valid = (|AlignerPlugin_logic_extractors_0_slicesOh);
    if(when_AlignerPlugin_l160) begin
      AlignerPlugin_logic_extractors_0_valid = 1'b0;
    end
    if(when_AlignerPlugin_l240) begin
      if(when_AlignerPlugin_l241) begin
        AlignerPlugin_logic_extractors_0_valid = 1'b0;
      end
    end
  end

  assign when_AlignerPlugin_l160 = (AlignerPlugin_api_haltIt || (AlignerPlugin_api_singleFetch && (! AlignerPlugin_logic_extractors_0_first)));
  assign when_AlignerPlugin_l171 = (decode_ctrls_0_up_isFiring && 1'b1);
  assign AlignerPlugin_logic_feeder_lanes_0_valid = AlignerPlugin_logic_extractors_0_valid;
  assign decode_ctrls_0_up_LANE_SEL_0 = AlignerPlugin_logic_feeder_lanes_0_valid;
  always @(*) begin
    decode_ctrls_0_up_Decode_INSTRUCTION_0 = AlignerPlugin_logic_extractors_0_ctx_instruction;
    if(AlignerPlugin_logic_feeder_lanes_0_isRvc) begin
      decode_ctrls_0_up_Decode_INSTRUCTION_0 = AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst;
    end
  end

  always @(*) begin
    decode_ctrls_0_up_Decode_DECOMPRESSION_FAULT_0 = 1'b0;
    if(AlignerPlugin_logic_feeder_lanes_0_isRvc) begin
      decode_ctrls_0_up_Decode_DECOMPRESSION_FAULT_0 = AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_illegal;
    end
  end

  always @(*) begin
    decode_ctrls_0_up_Decode_INSTRUCTION_RAW_0 = AlignerPlugin_logic_extractors_0_ctx_instruction;
    if(AlignerPlugin_logic_feeder_lanes_0_isRvc) begin
      decode_ctrls_0_up_Decode_INSTRUCTION_RAW_0[31 : 16] = 16'h0;
    end
  end

  assign AlignerPlugin_logic_feeder_lanes_0_isRvc = (AlignerPlugin_logic_extractors_0_ctx_instruction[1 : 0] != 2'b11);
  always @(*) begin
    AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(switch_Rvc_l55)
      5'h0 : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{{{{{{2'b00,AlignerPlugin_logic_extractors_0_ctx_instruction[10 : 7]},AlignerPlugin_logic_extractors_0_ctx_instruction[12 : 11]},AlignerPlugin_logic_extractors_0_ctx_instruction[5]},AlignerPlugin_logic_extractors_0_ctx_instruction[6]},2'b00},5'h02},3'b000},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_1},7'h13};
      end
      5'h02 : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_2,_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst},3'b010},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_1},7'h03};
      end
      5'h03 : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_3,_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst},3'b011},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_1},7'h03};
      end
      5'h05 : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_3[11 : 5],_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_1},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst},3'b011},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_3[4 : 0]},7'h27};
      end
      5'h06 : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_2[11 : 5],_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_1},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst},3'b010},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_2[4 : 0]},7'h23};
      end
      5'h07 : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_3[11 : 5],_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_1},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst},3'b011},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_3[4 : 0]},7'h23};
      end
      5'h08 : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_5,AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7]},3'b000},AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7]},7'h13};
      end
      5'h09 : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_5,AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7]},3'b000},AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7]},7'h1b};
      end
      5'h0a : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_5,5'h0},3'b000},AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7]},7'h13};
      end
      5'h0b : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = ((AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7] == 5'h02) ? {{{{{{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_19,_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_20},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_21},AlignerPlugin_logic_extractors_0_ctx_instruction[6]},4'b0000},AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7]},3'b000},AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7]},7'h13} : {{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_22[31 : 12],AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7]},7'h37});
      end
      5'h0c : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_23;
      end
      5'h0d : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_12[20],_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_12[10 : 1]},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_12[11]},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_12[19 : 12]},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_16},7'h6f};
      end
      5'h0e : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_15[12],_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_15[10 : 5]},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_16},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst},3'b000},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_15[4 : 1]},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_15[11]},7'h63};
      end
      5'h0f : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_15[12],_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_15[10 : 5]},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_16},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst},3'b001},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_15[4 : 1]},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_15[11]},7'h63};
      end
      5'h10 : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{{{6'h0,AlignerPlugin_logic_extractors_0_ctx_instruction[12]},AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 2]},AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7]},3'b001},AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7]},7'h13};
      end
      5'h12 : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{{{{{4'b0000,AlignerPlugin_logic_extractors_0_ctx_instruction[3 : 2]},AlignerPlugin_logic_extractors_0_ctx_instruction[12]},AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 4]},2'b00},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_17},3'b010},AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7]},7'h03};
      end
      5'h13 : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{{{{{3'b000,AlignerPlugin_logic_extractors_0_ctx_instruction[4 : 2]},AlignerPlugin_logic_extractors_0_ctx_instruction[12]},AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 5]},3'b000},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_17},3'b011},AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7]},7'h03};
      end
      5'h14 : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = ((AlignerPlugin_logic_extractors_0_ctx_instruction[12 : 2] == 11'h400) ? 32'h00100073 : ((AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 2] == 5'h0) ? {{{{12'h0,AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7]},3'b000},(AlignerPlugin_logic_extractors_0_ctx_instruction[12] ? 5'h01 : _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_16)},7'h67} : {{{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_27,_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_28},(_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_29 ? _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_30 : _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_16)},3'b000},AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7]},7'h33}));
      end
      5'h16 : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_31[11 : 5],AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 2]},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_17},3'b010},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_32[4 : 0]},7'h23};
      end
      5'h17 : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_33[11 : 5],AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 2]},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_17},3'b011},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_34[4 : 0]},7'h23};
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_illegal = 1'b0;
    case(switch_Rvc_l55)
      5'h0 : begin
        if(when_Rvc_l59) begin
          AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_illegal = 1'b1;
        end
      end
      5'h02 : begin
      end
      5'h03 : begin
      end
      5'h05 : begin
      end
      5'h06 : begin
      end
      5'h07 : begin
      end
      5'h08 : begin
      end
      5'h09 : begin
        if(when_Rvc_l73) begin
          AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_illegal = 1'b1;
        end
      end
      5'h0a : begin
      end
      5'h0b : begin
        if(when_Rvc_l80) begin
          AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_illegal = 1'b1;
        end
      end
      5'h0c : begin
      end
      5'h0d : begin
      end
      5'h0e : begin
      end
      5'h0f : begin
      end
      5'h10 : begin
      end
      5'h12 : begin
        if(when_Rvc_l101) begin
          AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_illegal = 1'b1;
        end
      end
      5'h13 : begin
        if(when_Rvc_l106) begin
          AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_illegal = 1'b1;
        end
      end
      5'h14 : begin
        if(when_Rvc_l114) begin
          AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_illegal = 1'b1;
        end
      end
      5'h16 : begin
      end
      5'h17 : begin
      end
      default : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_illegal = 1'b1;
      end
    endcase
  end

  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {2'b01,AlignerPlugin_logic_extractors_0_ctx_instruction[9 : 7]};
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_1 = {2'b01,AlignerPlugin_logic_extractors_0_ctx_instruction[4 : 2]};
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_2 = {{{{5'h0,AlignerPlugin_logic_extractors_0_ctx_instruction[5]},AlignerPlugin_logic_extractors_0_ctx_instruction[12 : 10]},AlignerPlugin_logic_extractors_0_ctx_instruction[6]},2'b00};
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_3 = {{{4'b0000,AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 5]},AlignerPlugin_logic_extractors_0_ctx_instruction[12 : 10]},3'b000};
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_4 = AlignerPlugin_logic_extractors_0_ctx_instruction[12];
  always @(*) begin
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_5[11] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_4;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_5[10] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_4;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_5[9] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_4;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_5[8] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_4;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_5[7] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_4;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_5[6] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_4;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_5[5] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_4;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_5[4 : 0] = AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 2];
  end

  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_6 = AlignerPlugin_logic_extractors_0_ctx_instruction[12];
  always @(*) begin
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_7[14] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_7[13] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_7[12] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_7[11] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_7[10] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_7[9] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_7[8] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_7[7] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_7[6] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_7[5] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_7[4] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_7[3] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_7[2] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_7[1] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_7[0] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_6;
  end

  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_8 = AlignerPlugin_logic_extractors_0_ctx_instruction[12];
  always @(*) begin
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_9[2] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_8;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_9[1] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_8;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_9[0] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_8;
  end

  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10 = AlignerPlugin_logic_extractors_0_ctx_instruction[12];
  always @(*) begin
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_11[9] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_11[8] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_11[7] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_11[6] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_11[5] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_11[4] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_11[3] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_11[2] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_11[1] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_11[0] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10;
  end

  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_12 = {{{{{{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_11,AlignerPlugin_logic_extractors_0_ctx_instruction[8]},AlignerPlugin_logic_extractors_0_ctx_instruction[10 : 9]},AlignerPlugin_logic_extractors_0_ctx_instruction[6]},AlignerPlugin_logic_extractors_0_ctx_instruction[7]},AlignerPlugin_logic_extractors_0_ctx_instruction[2]},AlignerPlugin_logic_extractors_0_ctx_instruction[11]},AlignerPlugin_logic_extractors_0_ctx_instruction[5 : 3]},1'b0};
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_13 = AlignerPlugin_logic_extractors_0_ctx_instruction[12];
  always @(*) begin
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_14[4] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_13;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_14[3] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_13;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_14[2] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_13;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_14[1] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_13;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_14[0] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_13;
  end

  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_15 = {{{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_14,AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 5]},AlignerPlugin_logic_extractors_0_ctx_instruction[2]},AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 10]},AlignerPlugin_logic_extractors_0_ctx_instruction[4 : 3]},1'b0};
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_16 = 5'h0;
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_17 = 5'h02;
  assign switch_Rvc_l55 = {AlignerPlugin_logic_extractors_0_ctx_instruction[1 : 0],AlignerPlugin_logic_extractors_0_ctx_instruction[15 : 13]};
  assign when_Rvc_l59 = (AlignerPlugin_logic_extractors_0_ctx_instruction[12 : 5] == 8'h0);
  assign when_Rvc_l73 = (AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7] == 5'h0);
  assign when_Rvc_l80 = ((AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 2] == 5'h0) && (AlignerPlugin_logic_extractors_0_ctx_instruction[12] == 1'b0));
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_18 = {{{{_zz__zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_18,_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst},3'b101},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst},7'h13};
  assign when_Rvc_l101 = (AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7] == 5'h0);
  assign when_Rvc_l106 = (AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7] == 5'h0);
  assign when_Rvc_l114 = (((AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7] == 5'h0) && (AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 2] == 5'h0)) && (AlignerPlugin_logic_extractors_0_ctx_instruction[12] == 1'b0));
  assign _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0 = AlignerPlugin_logic_extractors_0_localMask;
  assign _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_1 = {_zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0[0],_zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0[1]};
  assign _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_2 = _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_1[0];
  always @(*) begin
    _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_3[0] = (_zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_2 && (! 1'b0));
    _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_3[1] = (_zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_1[1] && (! _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_2));
  end

  assign _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_4 = _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_3;
  assign _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_5 = _zz__zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_5[1];
  assign decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0 = _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_5;
  assign decode_ctrls_0_up_PC_0 = AlignerPlugin_logic_extractors_0_ctx_pc;
  assign decode_ctrls_0_up_Decode_DOP_ID_0 = AlignerPlugin_logic_feeder_harts_0_dopId;
  assign decode_ctrls_0_up_Fetch_ID_0 = AlignerPlugin_logic_extractors_0_ctx_hm_Fetch_ID;
  assign decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_0_0 = AlignerPlugin_logic_extractors_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_0;
  assign decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_0_1 = AlignerPlugin_logic_extractors_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_1;
  assign decode_ctrls_0_up_Prediction_BRANCH_HISTORY_0 = AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_BRANCH_HISTORY;
  assign decode_ctrls_0_up_Prediction_WORD_SLICES_BRANCH_0 = AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_SLICES_BRANCH;
  assign decode_ctrls_0_up_Prediction_WORD_SLICES_TAKEN_0 = AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_SLICES_TAKEN;
  assign decode_ctrls_0_up_Prediction_WORD_JUMP_PC_0 = AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_JUMP_PC;
  assign decode_ctrls_0_up_Prediction_WORD_JUMPED_0 = AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_JUMPED;
  assign decode_ctrls_0_up_Prediction_WORD_JUMP_SLICE_0 = AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_JUMP_SLICE;
  assign decode_ctrls_0_up_TRAP_0 = AlignerPlugin_logic_extractors_0_ctx_trap;
  assign AlignerPlugin_logic_feeder_lanes_0_onBtb_pcLastSlice = (decode_ctrls_0_up_PC_0[1 : 1] + decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0);
  assign AlignerPlugin_logic_feeder_lanes_0_onBtb_didPrediction = (decode_ctrls_0_up_Prediction_WORD_JUMP_SLICE_0 <= AlignerPlugin_logic_feeder_lanes_0_onBtb_pcLastSlice);
  assign decode_ctrls_0_up_Prediction_ALIGNED_JUMPED_0 = (decode_ctrls_0_up_Prediction_WORD_JUMPED_0 && AlignerPlugin_logic_feeder_lanes_0_onBtb_didPrediction);
  assign decode_ctrls_0_up_Prediction_ALIGNED_JUMPED_PC_0 = decode_ctrls_0_up_Prediction_WORD_JUMP_PC_0;
  assign decode_ctrls_0_up_Prediction_ALIGNED_SLICES_BRANCH_0 = decode_ctrls_0_up_Prediction_WORD_SLICES_BRANCH_0;
  assign decode_ctrls_0_up_Prediction_ALIGNED_SLICES_TAKEN_0 = decode_ctrls_0_up_Prediction_WORD_SLICES_TAKEN_0;
  assign decode_ctrls_0_up_Prediction_ALIGN_REDO_0 = AlignerPlugin_logic_extractors_0_redo;
  assign decode_ctrls_0_up_valid = (|AlignerPlugin_logic_feeder_lanes_0_valid);
  assign _zz_AlignerPlugin_logic_slices_data_0 = {fetch_logic_ctrls_2_down_Fetch_WORD,AlignerPlugin_logic_buffer_data};
  assign AlignerPlugin_logic_slices_data_0 = _zz_AlignerPlugin_logic_slices_data_0[15 : 0];
  assign AlignerPlugin_logic_slices_data_1 = _zz_AlignerPlugin_logic_slices_data_0[31 : 16];
  assign AlignerPlugin_logic_slices_data_2 = _zz_AlignerPlugin_logic_slices_data_0[47 : 32];
  assign AlignerPlugin_logic_slices_data_3 = _zz_AlignerPlugin_logic_slices_data_0[63 : 48];
  assign AlignerPlugin_logic_slices_mask = {(fetch_logic_ctrls_2_down_isValid ? fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK : 2'b00),AlignerPlugin_logic_buffer_mask};
  assign AlignerPlugin_logic_slices_last = {fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_LAST,AlignerPlugin_logic_buffer_last};
  assign when_AlignerPlugin_l240 = (! fetch_logic_ctrls_2_down_valid);
  assign when_AlignerPlugin_l241 = (AlignerPlugin_logic_extractors_0_usageMask[3 : 2] != 2'b00);
  assign AlignerPlugin_logic_buffer_downFire = (decode_ctrls_0_up_isReady || decode_ctrls_0_up_isCancel);
  assign AlignerPlugin_logic_buffer_usedMask = (AlignerPlugin_logic_extractors_0_valid ? AlignerPlugin_logic_extractors_0_usageMask : 4'b0000);
  assign AlignerPlugin_logic_buffer_haltUp = ((|(AlignerPlugin_logic_buffer_mask & (~ (AlignerPlugin_logic_buffer_downFire ? AlignerPlugin_logic_buffer_usedMask[1 : 0] : 2'b00)))) || AlignerPlugin_api_haltIt);
  assign fetch_logic_ctrls_2_down_ready = ((! fetch_logic_ctrls_2_down_valid) || (! AlignerPlugin_logic_buffer_haltUp));
  assign when_AlignerPlugin_l256 = ((fetch_logic_ctrls_2_down_isValid && fetch_logic_ctrls_2_down_isReady) && (! fetch_logic_ctrls_2_down_isCancel));
  assign early0_EnvPlugin_logic_trapPort_payload_tval = (((execute_ctrl2_down_early0_EnvPlugin_OP_lane0 == EnvPluginOp_EBREAK) ? execute_ctrl2_down_PC_lane0 : 39'h0) | _zz_early0_EnvPlugin_logic_trapPort_payload_tval);
  always @(*) begin
    early0_EnvPlugin_logic_trapPort_payload_code = 4'b0010;
    case(execute_ctrl2_down_early0_EnvPlugin_OP_lane0)
      EnvPluginOp_EBREAK : begin
        early0_EnvPlugin_logic_trapPort_payload_code = 4'b0011;
      end
      EnvPluginOp_ECALL : begin
        early0_EnvPlugin_logic_trapPort_payload_code = (_zz_early0_EnvPlugin_logic_trapPort_payload_code | 4'b1000);
      end
      EnvPluginOp_PRIV_RET : begin
        if(when_EnvPlugin_l86) begin
          early0_EnvPlugin_logic_trapPort_payload_code = 4'b0001;
        end
      end
      EnvPluginOp_WFI : begin
        if(when_EnvPlugin_l95) begin
          early0_EnvPlugin_logic_trapPort_payload_code = 4'b1000;
        end
      end
      EnvPluginOp_FENCE_I : begin
        early0_EnvPlugin_logic_trapPort_payload_code = 4'b0010;
      end
      default : begin
        if(when_EnvPlugin_l110) begin
          early0_EnvPlugin_logic_trapPort_payload_code = 4'b0110;
        end
      end
    endcase
  end

  always @(*) begin
    early0_EnvPlugin_logic_trapPort_payload_arg = 3'bxxx;
    case(execute_ctrl2_down_early0_EnvPlugin_OP_lane0)
      EnvPluginOp_EBREAK : begin
      end
      EnvPluginOp_ECALL : begin
      end
      EnvPluginOp_PRIV_RET : begin
        if(when_EnvPlugin_l86) begin
          early0_EnvPlugin_logic_trapPort_payload_arg[1 : 0] = early0_EnvPlugin_logic_exe_xretPriv;
        end
      end
      EnvPluginOp_WFI : begin
      end
      EnvPluginOp_FENCE_I : begin
      end
      default : begin
      end
    endcase
  end

  assign early0_EnvPlugin_logic_exe_privilege = PrivilegedPlugin_logic_harts_0_privilege;
  assign early0_EnvPlugin_logic_exe_xretPriv = execute_ctrl2_down_Decode_UOP_lane0[29 : 28];
  always @(*) begin
    early0_EnvPlugin_logic_exe_commit = 1'b0;
    case(execute_ctrl2_down_early0_EnvPlugin_OP_lane0)
      EnvPluginOp_EBREAK : begin
      end
      EnvPluginOp_ECALL : begin
      end
      EnvPluginOp_PRIV_RET : begin
        if(when_EnvPlugin_l86) begin
          early0_EnvPlugin_logic_exe_commit = 1'b1;
        end
      end
      EnvPluginOp_WFI : begin
        if(when_EnvPlugin_l95) begin
          early0_EnvPlugin_logic_exe_commit = 1'b1;
        end
      end
      EnvPluginOp_FENCE_I : begin
        early0_EnvPlugin_logic_exe_commit = 1'b1;
      end
      default : begin
        if(when_EnvPlugin_l110) begin
          early0_EnvPlugin_logic_exe_commit = 1'b1;
        end
      end
    endcase
  end

  assign early0_EnvPlugin_logic_exe_retKo = ((PrivilegedPlugin_logic_harts_0_m_status_tsr && (early0_EnvPlugin_logic_exe_privilege == 2'b01)) && (early0_EnvPlugin_logic_exe_xretPriv == 2'b01));
  assign early0_EnvPlugin_logic_exe_vmaKo = (((early0_EnvPlugin_logic_exe_privilege == 2'b01) && PrivilegedPlugin_logic_harts_0_m_status_tvm) || (early0_EnvPlugin_logic_exe_privilege == 2'b00));
  assign when_EnvPlugin_l86 = ((early0_EnvPlugin_logic_exe_xretPriv <= PrivilegedPlugin_logic_harts_0_privilege) && (! early0_EnvPlugin_logic_exe_retKo));
  assign when_EnvPlugin_l95 = ((early0_EnvPlugin_logic_exe_privilege == 2'b11) || ((! PrivilegedPlugin_logic_harts_0_m_status_tw) && (1'b0 || (early0_EnvPlugin_logic_exe_privilege == 2'b01))));
  assign when_EnvPlugin_l110 = (! early0_EnvPlugin_logic_exe_vmaKo);
  assign when_EnvPlugin_l119 = (execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_down_early0_EnvPlugin_SEL_lane0);
  assign when_EnvPlugin_l123 = (! early0_EnvPlugin_logic_exe_commit);
  assign PmpPlugin_logic_isMachine = (PrivilegedPlugin_logic_harts_0_privilege == 2'b11);
  assign PmpPlugin_logic_instructionShouldHit = (! PmpPlugin_logic_isMachine);
  assign PmpPlugin_logic_dataShouldHit = ((! PmpPlugin_logic_isMachine) || (PrivilegedPlugin_logic_harts_0_m_status_mprv && (PrivilegedPlugin_logic_harts_0_m_status_mpp != 2'b11)));
  assign FetchL1Plugin_logic_pmpPort_logic_dataShouldHitPort = (PmpPlugin_logic_dataShouldHit || 1'b0);
  assign FetchL1Plugin_logic_pmpPort_logic_torCmpAddress = (fetch_logic_ctrls_1_down_MMU_TRANSLATED >>> 4'd12);
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_napot_MATCH = ((_zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_napot_MATCH[31 : 12] ^ fetch_logic_ctrls_1_down_MMU_TRANSLATED[31 : 12]) & PmpPlugin_logic_entries_0_mask);
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_napot_HIT = (fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_napot_MATCH == 20'h0);
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_tor_BIGGER = (FetchL1Plugin_logic_pmpPort_logic_torCmpAddress < _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_tor_BIGGER);
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_tor_HIT = (fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_tor_BIGGER && 1'b1);
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_HIT_ANY = ((PmpPlugin_logic_entries_0_isNapot && fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_napot_HIT) || (PmpPlugin_logic_entries_0_isTor && fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_tor_HIT));
  assign FetchL1Plugin_logic_pmpPort_logic_onEntries_0_instructionCheck = (PmpPlugin_logic_entries_0_cfg_locked || PmpPlugin_logic_instructionShouldHit);
  assign FetchL1Plugin_logic_pmpPort_logic_onEntries_0_dataCheck = (PmpPlugin_logic_entries_0_cfg_locked || FetchL1Plugin_logic_pmpPort_logic_dataShouldHitPort);
  assign FetchL1Plugin_logic_pmpPort_logic_onEntries_0_normalRwx = ((((! 1'b1) || PmpPlugin_logic_entries_0_cfg_execute) || (! FetchL1Plugin_logic_pmpPort_logic_onEntries_0_instructionCheck)) && ((((! 1'b0) || PmpPlugin_logic_entries_0_cfg_write) && ((! 1'b0) || PmpPlugin_logic_entries_0_cfg_read)) || (! FetchL1Plugin_logic_pmpPort_logic_onEntries_0_dataCheck)));
  assign fetch_logic_ctrls_0_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_PERM_OK = FetchL1Plugin_logic_pmpPort_logic_onEntries_0_normalRwx;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_napot_MATCH = ((_zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_napot_MATCH[31 : 12] ^ fetch_logic_ctrls_1_down_MMU_TRANSLATED[31 : 12]) & PmpPlugin_logic_entries_1_mask);
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_napot_HIT = (fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_napot_MATCH == 20'h0);
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_tor_BIGGER = (FetchL1Plugin_logic_pmpPort_logic_torCmpAddress < _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_tor_BIGGER);
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_tor_HIT = (fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_tor_BIGGER && (! fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_tor_BIGGER));
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_HIT_ANY = ((PmpPlugin_logic_entries_1_isNapot && fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_napot_HIT) || (PmpPlugin_logic_entries_1_isTor && fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_tor_HIT));
  assign FetchL1Plugin_logic_pmpPort_logic_onEntries_1_instructionCheck = (PmpPlugin_logic_entries_1_cfg_locked || PmpPlugin_logic_instructionShouldHit);
  assign FetchL1Plugin_logic_pmpPort_logic_onEntries_1_dataCheck = (PmpPlugin_logic_entries_1_cfg_locked || FetchL1Plugin_logic_pmpPort_logic_dataShouldHitPort);
  assign FetchL1Plugin_logic_pmpPort_logic_onEntries_1_normalRwx = ((((! 1'b1) || PmpPlugin_logic_entries_1_cfg_execute) || (! FetchL1Plugin_logic_pmpPort_logic_onEntries_1_instructionCheck)) && ((((! 1'b0) || PmpPlugin_logic_entries_1_cfg_write) && ((! 1'b0) || PmpPlugin_logic_entries_1_cfg_read)) || (! FetchL1Plugin_logic_pmpPort_logic_onEntries_1_dataCheck)));
  assign fetch_logic_ctrls_0_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_PERM_OK = FetchL1Plugin_logic_pmpPort_logic_onEntries_1_normalRwx;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_napot_MATCH = ((_zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_napot_MATCH[31 : 12] ^ fetch_logic_ctrls_1_down_MMU_TRANSLATED[31 : 12]) & PmpPlugin_logic_entries_2_mask);
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_napot_HIT = (fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_napot_MATCH == 20'h0);
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_tor_BIGGER = (FetchL1Plugin_logic_pmpPort_logic_torCmpAddress < _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_tor_BIGGER);
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_tor_HIT = (fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_tor_BIGGER && (! fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_tor_BIGGER));
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_HIT_ANY = ((PmpPlugin_logic_entries_2_isNapot && fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_napot_HIT) || (PmpPlugin_logic_entries_2_isTor && fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_tor_HIT));
  assign FetchL1Plugin_logic_pmpPort_logic_onEntries_2_instructionCheck = (PmpPlugin_logic_entries_2_cfg_locked || PmpPlugin_logic_instructionShouldHit);
  assign FetchL1Plugin_logic_pmpPort_logic_onEntries_2_dataCheck = (PmpPlugin_logic_entries_2_cfg_locked || FetchL1Plugin_logic_pmpPort_logic_dataShouldHitPort);
  assign FetchL1Plugin_logic_pmpPort_logic_onEntries_2_normalRwx = ((((! 1'b1) || PmpPlugin_logic_entries_2_cfg_execute) || (! FetchL1Plugin_logic_pmpPort_logic_onEntries_2_instructionCheck)) && ((((! 1'b0) || PmpPlugin_logic_entries_2_cfg_write) && ((! 1'b0) || PmpPlugin_logic_entries_2_cfg_read)) || (! FetchL1Plugin_logic_pmpPort_logic_onEntries_2_dataCheck)));
  assign fetch_logic_ctrls_0_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_PERM_OK = FetchL1Plugin_logic_pmpPort_logic_onEntries_2_normalRwx;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_napot_MATCH = ((_zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_napot_MATCH[31 : 12] ^ fetch_logic_ctrls_1_down_MMU_TRANSLATED[31 : 12]) & PmpPlugin_logic_entries_3_mask);
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_napot_HIT = (fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_napot_MATCH == 20'h0);
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_tor_BIGGER = (FetchL1Plugin_logic_pmpPort_logic_torCmpAddress < _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_tor_BIGGER);
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_tor_HIT = (fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_tor_BIGGER && (! fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_tor_BIGGER));
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_HIT_ANY = ((PmpPlugin_logic_entries_3_isNapot && fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_napot_HIT) || (PmpPlugin_logic_entries_3_isTor && fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_tor_HIT));
  assign FetchL1Plugin_logic_pmpPort_logic_onEntries_3_instructionCheck = (PmpPlugin_logic_entries_3_cfg_locked || PmpPlugin_logic_instructionShouldHit);
  assign FetchL1Plugin_logic_pmpPort_logic_onEntries_3_dataCheck = (PmpPlugin_logic_entries_3_cfg_locked || FetchL1Plugin_logic_pmpPort_logic_dataShouldHitPort);
  assign FetchL1Plugin_logic_pmpPort_logic_onEntries_3_normalRwx = ((((! 1'b1) || PmpPlugin_logic_entries_3_cfg_execute) || (! FetchL1Plugin_logic_pmpPort_logic_onEntries_3_instructionCheck)) && ((((! 1'b0) || PmpPlugin_logic_entries_3_cfg_write) && ((! 1'b0) || PmpPlugin_logic_entries_3_cfg_read)) || (! FetchL1Plugin_logic_pmpPort_logic_onEntries_3_dataCheck)));
  assign fetch_logic_ctrls_0_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_PERM_OK = FetchL1Plugin_logic_pmpPort_logic_onEntries_3_normalRwx;
  assign fetch_logic_ctrls_0_down_FetchL1Plugin_logic_pmpPort_logic_NEED_HIT = ((PmpPlugin_logic_instructionShouldHit && 1'b1) || (FetchL1Plugin_logic_pmpPort_logic_dataShouldHitPort && (1'b0 || 1'b0)));
  assign FetchL1Plugin_logic_pmpPort_logic_onCtrl_hits = {fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_HIT_ANY,{fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_HIT_ANY,{fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_HIT_ANY,fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_HIT_ANY}}};
  assign _zz_FetchL1Plugin_logic_pmpPort_logic_onCtrl_hits_bools_0 = FetchL1Plugin_logic_pmpPort_logic_onCtrl_hits;
  assign FetchL1Plugin_logic_pmpPort_logic_onCtrl_hits_bools_0 = _zz_FetchL1Plugin_logic_pmpPort_logic_onCtrl_hits_bools_0[0];
  assign FetchL1Plugin_logic_pmpPort_logic_onCtrl_hits_bools_1 = _zz_FetchL1Plugin_logic_pmpPort_logic_onCtrl_hits_bools_0[1];
  assign FetchL1Plugin_logic_pmpPort_logic_onCtrl_hits_bools_2 = _zz_FetchL1Plugin_logic_pmpPort_logic_onCtrl_hits_bools_0[2];
  assign FetchL1Plugin_logic_pmpPort_logic_onCtrl_hits_bools_3 = _zz_FetchL1Plugin_logic_pmpPort_logic_onCtrl_hits_bools_0[3];
  always @(*) begin
    _zz_FetchL1Plugin_logic_pmpPort_logic_onCtrl_oh[0] = (FetchL1Plugin_logic_pmpPort_logic_onCtrl_hits_bools_0 && (! 1'b0));
    _zz_FetchL1Plugin_logic_pmpPort_logic_onCtrl_oh[1] = (FetchL1Plugin_logic_pmpPort_logic_onCtrl_hits_bools_1 && (! FetchL1Plugin_logic_pmpPort_logic_onCtrl_hits_bools_0));
    _zz_FetchL1Plugin_logic_pmpPort_logic_onCtrl_oh[2] = (FetchL1Plugin_logic_pmpPort_logic_onCtrl_hits_bools_2 && (! FetchL1Plugin_logic_pmpPort_logic_onCtrl_hits_range_0_to_1));
    _zz_FetchL1Plugin_logic_pmpPort_logic_onCtrl_oh[3] = (FetchL1Plugin_logic_pmpPort_logic_onCtrl_hits_bools_3 && (! FetchL1Plugin_logic_pmpPort_logic_onCtrl_hits_range_0_to_2));
  end

  assign FetchL1Plugin_logic_pmpPort_logic_onCtrl_hits_range_0_to_1 = (|{FetchL1Plugin_logic_pmpPort_logic_onCtrl_hits_bools_1,FetchL1Plugin_logic_pmpPort_logic_onCtrl_hits_bools_0});
  assign FetchL1Plugin_logic_pmpPort_logic_onCtrl_hits_range_0_to_2 = (|{FetchL1Plugin_logic_pmpPort_logic_onCtrl_hits_bools_2,{FetchL1Plugin_logic_pmpPort_logic_onCtrl_hits_bools_1,FetchL1Plugin_logic_pmpPort_logic_onCtrl_hits_bools_0}});
  assign FetchL1Plugin_logic_pmpPort_logic_onCtrl_oh = _zz_FetchL1Plugin_logic_pmpPort_logic_onCtrl_oh;
  assign _zz_fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_ACCESS_FAULT = FetchL1Plugin_logic_pmpPort_logic_onCtrl_oh[0];
  assign _zz_fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_ACCESS_FAULT_1 = FetchL1Plugin_logic_pmpPort_logic_onCtrl_oh[1];
  assign _zz_fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_ACCESS_FAULT_2 = FetchL1Plugin_logic_pmpPort_logic_onCtrl_oh[2];
  assign _zz_fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_ACCESS_FAULT_3 = FetchL1Plugin_logic_pmpPort_logic_onCtrl_oh[3];
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_ACCESS_FAULT = ((fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_NEED_HIT || _zz_fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_ACCESS_FAULT_4[0]) && (! _zz_fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_ACCESS_FAULT_5[0]));
  assign LsuPlugin_logic_pmpPort_logic_dataShouldHitPort = (PmpPlugin_logic_dataShouldHit || execute_ctrl2_down_LsuPlugin_logic_FROM_ACCESS_lane0);
  assign LsuPlugin_logic_pmpPort_logic_torCmpAddress = (execute_ctrl3_down_MMU_TRANSLATED_lane0 >>> 4'd12);
  assign execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_0_napot_MATCH_lane0 = ((_zz_execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_0_napot_MATCH_lane0[31 : 12] ^ execute_ctrl3_down_MMU_TRANSLATED_lane0[31 : 12]) & PmpPlugin_logic_entries_0_mask);
  assign execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_0_napot_HIT_lane0 = (execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_0_napot_MATCH_lane0 == 20'h0);
  assign execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_0_tor_BIGGER_lane0 = (LsuPlugin_logic_pmpPort_logic_torCmpAddress < _zz_execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_0_tor_BIGGER_lane0);
  assign execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_0_tor_HIT_lane0 = (execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_0_tor_BIGGER_lane0 && 1'b1);
  assign execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_0_HIT_ANY_lane0 = ((PmpPlugin_logic_entries_0_isNapot && execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_0_napot_HIT_lane0) || (PmpPlugin_logic_entries_0_isTor && execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_0_tor_HIT_lane0));
  assign LsuPlugin_logic_pmpPort_logic_onEntries_0_instructionCheck = (PmpPlugin_logic_entries_0_cfg_locked || PmpPlugin_logic_instructionShouldHit);
  assign LsuPlugin_logic_pmpPort_logic_onEntries_0_dataCheck = (PmpPlugin_logic_entries_0_cfg_locked || LsuPlugin_logic_pmpPort_logic_dataShouldHitPort);
  assign LsuPlugin_logic_pmpPort_logic_onEntries_0_normalRwx = ((((! 1'b0) || PmpPlugin_logic_entries_0_cfg_execute) || (! LsuPlugin_logic_pmpPort_logic_onEntries_0_instructionCheck)) && ((((! execute_ctrl2_down_LsuL1_STORE_lane0) || PmpPlugin_logic_entries_0_cfg_write) && ((! execute_ctrl2_down_LsuL1_LOAD_lane0) || PmpPlugin_logic_entries_0_cfg_read)) || (! LsuPlugin_logic_pmpPort_logic_onEntries_0_dataCheck)));
  assign execute_ctrl2_down_LsuPlugin_logic_pmpPort_logic_onEntries_0_PERM_OK_lane0 = LsuPlugin_logic_pmpPort_logic_onEntries_0_normalRwx;
  assign execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_1_napot_MATCH_lane0 = ((_zz_execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_1_napot_MATCH_lane0[31 : 12] ^ execute_ctrl3_down_MMU_TRANSLATED_lane0[31 : 12]) & PmpPlugin_logic_entries_1_mask);
  assign execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_1_napot_HIT_lane0 = (execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_1_napot_MATCH_lane0 == 20'h0);
  assign execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_1_tor_BIGGER_lane0 = (LsuPlugin_logic_pmpPort_logic_torCmpAddress < _zz_execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_1_tor_BIGGER_lane0);
  assign execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_1_tor_HIT_lane0 = (execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_1_tor_BIGGER_lane0 && (! execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_0_tor_BIGGER_lane0));
  assign execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_1_HIT_ANY_lane0 = ((PmpPlugin_logic_entries_1_isNapot && execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_1_napot_HIT_lane0) || (PmpPlugin_logic_entries_1_isTor && execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_1_tor_HIT_lane0));
  assign LsuPlugin_logic_pmpPort_logic_onEntries_1_instructionCheck = (PmpPlugin_logic_entries_1_cfg_locked || PmpPlugin_logic_instructionShouldHit);
  assign LsuPlugin_logic_pmpPort_logic_onEntries_1_dataCheck = (PmpPlugin_logic_entries_1_cfg_locked || LsuPlugin_logic_pmpPort_logic_dataShouldHitPort);
  assign LsuPlugin_logic_pmpPort_logic_onEntries_1_normalRwx = ((((! 1'b0) || PmpPlugin_logic_entries_1_cfg_execute) || (! LsuPlugin_logic_pmpPort_logic_onEntries_1_instructionCheck)) && ((((! execute_ctrl2_down_LsuL1_STORE_lane0) || PmpPlugin_logic_entries_1_cfg_write) && ((! execute_ctrl2_down_LsuL1_LOAD_lane0) || PmpPlugin_logic_entries_1_cfg_read)) || (! LsuPlugin_logic_pmpPort_logic_onEntries_1_dataCheck)));
  assign execute_ctrl2_down_LsuPlugin_logic_pmpPort_logic_onEntries_1_PERM_OK_lane0 = LsuPlugin_logic_pmpPort_logic_onEntries_1_normalRwx;
  assign execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_2_napot_MATCH_lane0 = ((_zz_execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_2_napot_MATCH_lane0[31 : 12] ^ execute_ctrl3_down_MMU_TRANSLATED_lane0[31 : 12]) & PmpPlugin_logic_entries_2_mask);
  assign execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_2_napot_HIT_lane0 = (execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_2_napot_MATCH_lane0 == 20'h0);
  assign execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_2_tor_BIGGER_lane0 = (LsuPlugin_logic_pmpPort_logic_torCmpAddress < _zz_execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_2_tor_BIGGER_lane0);
  assign execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_2_tor_HIT_lane0 = (execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_2_tor_BIGGER_lane0 && (! execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_1_tor_BIGGER_lane0));
  assign execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_2_HIT_ANY_lane0 = ((PmpPlugin_logic_entries_2_isNapot && execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_2_napot_HIT_lane0) || (PmpPlugin_logic_entries_2_isTor && execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_2_tor_HIT_lane0));
  assign LsuPlugin_logic_pmpPort_logic_onEntries_2_instructionCheck = (PmpPlugin_logic_entries_2_cfg_locked || PmpPlugin_logic_instructionShouldHit);
  assign LsuPlugin_logic_pmpPort_logic_onEntries_2_dataCheck = (PmpPlugin_logic_entries_2_cfg_locked || LsuPlugin_logic_pmpPort_logic_dataShouldHitPort);
  assign LsuPlugin_logic_pmpPort_logic_onEntries_2_normalRwx = ((((! 1'b0) || PmpPlugin_logic_entries_2_cfg_execute) || (! LsuPlugin_logic_pmpPort_logic_onEntries_2_instructionCheck)) && ((((! execute_ctrl2_down_LsuL1_STORE_lane0) || PmpPlugin_logic_entries_2_cfg_write) && ((! execute_ctrl2_down_LsuL1_LOAD_lane0) || PmpPlugin_logic_entries_2_cfg_read)) || (! LsuPlugin_logic_pmpPort_logic_onEntries_2_dataCheck)));
  assign execute_ctrl2_down_LsuPlugin_logic_pmpPort_logic_onEntries_2_PERM_OK_lane0 = LsuPlugin_logic_pmpPort_logic_onEntries_2_normalRwx;
  assign execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_3_napot_MATCH_lane0 = ((_zz_execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_3_napot_MATCH_lane0[31 : 12] ^ execute_ctrl3_down_MMU_TRANSLATED_lane0[31 : 12]) & PmpPlugin_logic_entries_3_mask);
  assign execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_3_napot_HIT_lane0 = (execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_3_napot_MATCH_lane0 == 20'h0);
  assign execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_3_tor_BIGGER_lane0 = (LsuPlugin_logic_pmpPort_logic_torCmpAddress < _zz_execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_3_tor_BIGGER_lane0);
  assign execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_3_tor_HIT_lane0 = (execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_3_tor_BIGGER_lane0 && (! execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_2_tor_BIGGER_lane0));
  assign execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_3_HIT_ANY_lane0 = ((PmpPlugin_logic_entries_3_isNapot && execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_3_napot_HIT_lane0) || (PmpPlugin_logic_entries_3_isTor && execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_3_tor_HIT_lane0));
  assign LsuPlugin_logic_pmpPort_logic_onEntries_3_instructionCheck = (PmpPlugin_logic_entries_3_cfg_locked || PmpPlugin_logic_instructionShouldHit);
  assign LsuPlugin_logic_pmpPort_logic_onEntries_3_dataCheck = (PmpPlugin_logic_entries_3_cfg_locked || LsuPlugin_logic_pmpPort_logic_dataShouldHitPort);
  assign LsuPlugin_logic_pmpPort_logic_onEntries_3_normalRwx = ((((! 1'b0) || PmpPlugin_logic_entries_3_cfg_execute) || (! LsuPlugin_logic_pmpPort_logic_onEntries_3_instructionCheck)) && ((((! execute_ctrl2_down_LsuL1_STORE_lane0) || PmpPlugin_logic_entries_3_cfg_write) && ((! execute_ctrl2_down_LsuL1_LOAD_lane0) || PmpPlugin_logic_entries_3_cfg_read)) || (! LsuPlugin_logic_pmpPort_logic_onEntries_3_dataCheck)));
  assign execute_ctrl2_down_LsuPlugin_logic_pmpPort_logic_onEntries_3_PERM_OK_lane0 = LsuPlugin_logic_pmpPort_logic_onEntries_3_normalRwx;
  assign execute_ctrl2_down_LsuPlugin_logic_pmpPort_logic_NEED_HIT_lane0 = ((PmpPlugin_logic_instructionShouldHit && 1'b0) || (LsuPlugin_logic_pmpPort_logic_dataShouldHitPort && (execute_ctrl2_down_LsuL1_LOAD_lane0 || execute_ctrl2_down_LsuL1_STORE_lane0)));
  assign LsuPlugin_logic_pmpPort_logic_onCtrl_hits = {execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_3_HIT_ANY_lane0,{execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_2_HIT_ANY_lane0,{execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_1_HIT_ANY_lane0,execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_0_HIT_ANY_lane0}}};
  assign _zz_LsuPlugin_logic_pmpPort_logic_onCtrl_hits_bools_0 = LsuPlugin_logic_pmpPort_logic_onCtrl_hits;
  assign LsuPlugin_logic_pmpPort_logic_onCtrl_hits_bools_0 = _zz_LsuPlugin_logic_pmpPort_logic_onCtrl_hits_bools_0[0];
  assign LsuPlugin_logic_pmpPort_logic_onCtrl_hits_bools_1 = _zz_LsuPlugin_logic_pmpPort_logic_onCtrl_hits_bools_0[1];
  assign LsuPlugin_logic_pmpPort_logic_onCtrl_hits_bools_2 = _zz_LsuPlugin_logic_pmpPort_logic_onCtrl_hits_bools_0[2];
  assign LsuPlugin_logic_pmpPort_logic_onCtrl_hits_bools_3 = _zz_LsuPlugin_logic_pmpPort_logic_onCtrl_hits_bools_0[3];
  always @(*) begin
    _zz_LsuPlugin_logic_pmpPort_logic_onCtrl_oh[0] = (LsuPlugin_logic_pmpPort_logic_onCtrl_hits_bools_0 && (! 1'b0));
    _zz_LsuPlugin_logic_pmpPort_logic_onCtrl_oh[1] = (LsuPlugin_logic_pmpPort_logic_onCtrl_hits_bools_1 && (! LsuPlugin_logic_pmpPort_logic_onCtrl_hits_bools_0));
    _zz_LsuPlugin_logic_pmpPort_logic_onCtrl_oh[2] = (LsuPlugin_logic_pmpPort_logic_onCtrl_hits_bools_2 && (! LsuPlugin_logic_pmpPort_logic_onCtrl_hits_range_0_to_1));
    _zz_LsuPlugin_logic_pmpPort_logic_onCtrl_oh[3] = (LsuPlugin_logic_pmpPort_logic_onCtrl_hits_bools_3 && (! LsuPlugin_logic_pmpPort_logic_onCtrl_hits_range_0_to_2));
  end

  assign LsuPlugin_logic_pmpPort_logic_onCtrl_hits_range_0_to_1 = (|{LsuPlugin_logic_pmpPort_logic_onCtrl_hits_bools_1,LsuPlugin_logic_pmpPort_logic_onCtrl_hits_bools_0});
  assign LsuPlugin_logic_pmpPort_logic_onCtrl_hits_range_0_to_2 = (|{LsuPlugin_logic_pmpPort_logic_onCtrl_hits_bools_2,{LsuPlugin_logic_pmpPort_logic_onCtrl_hits_bools_1,LsuPlugin_logic_pmpPort_logic_onCtrl_hits_bools_0}});
  assign LsuPlugin_logic_pmpPort_logic_onCtrl_oh = _zz_LsuPlugin_logic_pmpPort_logic_onCtrl_oh;
  assign _zz_execute_ctrl4_down_LsuPlugin_logic_pmpPort_ACCESS_FAULT_lane0 = LsuPlugin_logic_pmpPort_logic_onCtrl_oh[0];
  assign _zz_execute_ctrl4_down_LsuPlugin_logic_pmpPort_ACCESS_FAULT_lane0_1 = LsuPlugin_logic_pmpPort_logic_onCtrl_oh[1];
  assign _zz_execute_ctrl4_down_LsuPlugin_logic_pmpPort_ACCESS_FAULT_lane0_2 = LsuPlugin_logic_pmpPort_logic_onCtrl_oh[2];
  assign _zz_execute_ctrl4_down_LsuPlugin_logic_pmpPort_ACCESS_FAULT_lane0_3 = LsuPlugin_logic_pmpPort_logic_onCtrl_oh[3];
  assign execute_ctrl4_down_LsuPlugin_logic_pmpPort_ACCESS_FAULT_lane0 = ((execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_NEED_HIT_lane0 || _zz_execute_ctrl4_down_LsuPlugin_logic_pmpPort_ACCESS_FAULT_lane0_4[0]) && (! _zz_execute_ctrl4_down_LsuPlugin_logic_pmpPort_ACCESS_FAULT_lane0_5[0]));
  assign LsuCachelessAxi4Plugin_logic_bridge_cmdHash = LsuPlugin_logic_bus_cmd_payload_address[10 : 3];
  assign LsuCachelessAxi4Plugin_logic_bridge_tracker_pendings_0_hazard = (LsuCachelessAxi4Plugin_logic_bridge_tracker_pendings_0_valid && (((LsuCachelessAxi4Plugin_logic_bridge_tracker_pendings_0_hash == LsuCachelessAxi4Plugin_logic_bridge_cmdHash) && (|(LsuCachelessAxi4Plugin_logic_bridge_tracker_pendings_0_mask & LsuPlugin_logic_bus_cmd_payload_mask))) || (LsuCachelessAxi4Plugin_logic_bridge_tracker_pendings_0_io && LsuPlugin_logic_bus_cmd_payload_io)));
  assign LsuCachelessAxi4Plugin_logic_bridge_tracker_hazard = (|LsuCachelessAxi4Plugin_logic_bridge_tracker_pendings_0_hazard);
  assign _zz_LsuPlugin_logic_bus_cmd_ready = (! LsuCachelessAxi4Plugin_logic_bridge_tracker_hazard);
  assign LsuPlugin_logic_bus_cmd_haltWhen_valid = (LsuPlugin_logic_bus_cmd_valid && _zz_LsuPlugin_logic_bus_cmd_ready);
  assign LsuPlugin_logic_bus_cmd_ready = (LsuPlugin_logic_bus_cmd_haltWhen_ready && _zz_LsuPlugin_logic_bus_cmd_ready);
  assign LsuPlugin_logic_bus_cmd_haltWhen_payload_write = LsuPlugin_logic_bus_cmd_payload_write;
  assign LsuPlugin_logic_bus_cmd_haltWhen_payload_address = LsuPlugin_logic_bus_cmd_payload_address;
  assign LsuPlugin_logic_bus_cmd_haltWhen_payload_data = LsuPlugin_logic_bus_cmd_payload_data;
  assign LsuPlugin_logic_bus_cmd_haltWhen_payload_size = LsuPlugin_logic_bus_cmd_payload_size;
  assign LsuPlugin_logic_bus_cmd_haltWhen_payload_mask = LsuPlugin_logic_bus_cmd_payload_mask;
  assign LsuPlugin_logic_bus_cmd_haltWhen_payload_io = LsuPlugin_logic_bus_cmd_payload_io;
  assign LsuPlugin_logic_bus_cmd_haltWhen_payload_fromHart = LsuPlugin_logic_bus_cmd_payload_fromHart;
  assign LsuPlugin_logic_bus_cmd_haltWhen_payload_uopId = LsuPlugin_logic_bus_cmd_payload_uopId;
  assign LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_valid = LsuPlugin_logic_bus_cmd_haltWhen_valid;
  assign LsuPlugin_logic_bus_cmd_haltWhen_ready = LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_ready;
  assign LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_payload_write = LsuPlugin_logic_bus_cmd_haltWhen_payload_write;
  assign LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_payload_address = LsuPlugin_logic_bus_cmd_haltWhen_payload_address;
  assign LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_payload_data = LsuPlugin_logic_bus_cmd_haltWhen_payload_data;
  assign LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_payload_size = LsuPlugin_logic_bus_cmd_haltWhen_payload_size;
  assign LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_payload_mask = LsuPlugin_logic_bus_cmd_haltWhen_payload_mask;
  assign LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_payload_io = LsuPlugin_logic_bus_cmd_haltWhen_payload_io;
  assign LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_payload_fromHart = LsuPlugin_logic_bus_cmd_haltWhen_payload_fromHart;
  assign LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_payload_uopId = LsuPlugin_logic_bus_cmd_haltWhen_payload_uopId;
  always @(*) begin
    LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_ready = 1'b1;
    if(when_Stream_l1253_2) begin
      LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_ready = 1'b0;
    end
    if(when_Stream_l1253_3) begin
      LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_ready = 1'b0;
    end
  end

  assign when_Stream_l1253_2 = ((! LsuCachelessAxi4Plugin_logic_bridge_cmdFork_ready) && LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_fork2_logic_linkEnable_0);
  assign when_Stream_l1253_3 = ((! LsuCachelessAxi4Plugin_logic_bridge_dataFork_ready) && LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_fork2_logic_linkEnable_1);
  assign LsuCachelessAxi4Plugin_logic_bridge_cmdFork_valid = (LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_valid && LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_fork2_logic_linkEnable_0);
  assign LsuCachelessAxi4Plugin_logic_bridge_cmdFork_payload_write = LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_payload_write;
  assign LsuCachelessAxi4Plugin_logic_bridge_cmdFork_payload_address = LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_payload_address;
  assign LsuCachelessAxi4Plugin_logic_bridge_cmdFork_payload_data = LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_payload_data;
  assign LsuCachelessAxi4Plugin_logic_bridge_cmdFork_payload_size = LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_payload_size;
  assign LsuCachelessAxi4Plugin_logic_bridge_cmdFork_payload_mask = LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_payload_mask;
  assign LsuCachelessAxi4Plugin_logic_bridge_cmdFork_payload_io = LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_payload_io;
  assign LsuCachelessAxi4Plugin_logic_bridge_cmdFork_payload_fromHart = LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_payload_fromHart;
  assign LsuCachelessAxi4Plugin_logic_bridge_cmdFork_payload_uopId = LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_payload_uopId;
  assign LsuCachelessAxi4Plugin_logic_bridge_cmdFork_fire = (LsuCachelessAxi4Plugin_logic_bridge_cmdFork_valid && LsuCachelessAxi4Plugin_logic_bridge_cmdFork_ready);
  assign LsuCachelessAxi4Plugin_logic_bridge_dataFork_valid = (LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_valid && LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_fork2_logic_linkEnable_1);
  assign LsuCachelessAxi4Plugin_logic_bridge_dataFork_payload_write = LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_payload_write;
  assign LsuCachelessAxi4Plugin_logic_bridge_dataFork_payload_address = LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_payload_address;
  assign LsuCachelessAxi4Plugin_logic_bridge_dataFork_payload_data = LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_payload_data;
  assign LsuCachelessAxi4Plugin_logic_bridge_dataFork_payload_size = LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_payload_size;
  assign LsuCachelessAxi4Plugin_logic_bridge_dataFork_payload_mask = LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_payload_mask;
  assign LsuCachelessAxi4Plugin_logic_bridge_dataFork_payload_io = LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_payload_io;
  assign LsuCachelessAxi4Plugin_logic_bridge_dataFork_payload_fromHart = LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_payload_fromHart;
  assign LsuCachelessAxi4Plugin_logic_bridge_dataFork_payload_uopId = LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_payload_uopId;
  assign LsuCachelessAxi4Plugin_logic_bridge_dataFork_fire = (LsuCachelessAxi4Plugin_logic_bridge_dataFork_valid && LsuCachelessAxi4Plugin_logic_bridge_dataFork_ready);
  assign LsuCachelessAxi4Plugin_logic_bridge_down_arw_valid = LsuCachelessAxi4Plugin_logic_bridge_cmdFork_valid;
  assign LsuCachelessAxi4Plugin_logic_bridge_cmdFork_ready = LsuCachelessAxi4Plugin_logic_bridge_down_arw_ready;
  assign LsuCachelessAxi4Plugin_logic_bridge_down_arw_payload_write = LsuCachelessAxi4Plugin_logic_bridge_cmdFork_payload_write;
  assign LsuCachelessAxi4Plugin_logic_bridge_down_arw_payload_prot = 3'b010;
  assign LsuCachelessAxi4Plugin_logic_bridge_down_arw_payload_cache = (LsuCachelessAxi4Plugin_logic_bridge_cmdFork_payload_io ? 4'b0000 : 4'b1111);
  assign LsuCachelessAxi4Plugin_logic_bridge_down_arw_payload_size = {1'd0, LsuCachelessAxi4Plugin_logic_bridge_cmdFork_payload_size};
  assign LsuCachelessAxi4Plugin_logic_bridge_down_arw_payload_addr = LsuCachelessAxi4Plugin_logic_bridge_cmdFork_payload_address;
  assign when_Stream_l581_1 = (! LsuCachelessAxi4Plugin_logic_bridge_dataFork_payload_write);
  always @(*) begin
    LsuCachelessAxi4Plugin_logic_bridge_dataStage_valid = LsuCachelessAxi4Plugin_logic_bridge_dataFork_valid;
    if(when_Stream_l581_1) begin
      LsuCachelessAxi4Plugin_logic_bridge_dataStage_valid = 1'b0;
    end
  end

  always @(*) begin
    LsuCachelessAxi4Plugin_logic_bridge_dataFork_ready = LsuCachelessAxi4Plugin_logic_bridge_dataStage_ready;
    if(when_Stream_l581_1) begin
      LsuCachelessAxi4Plugin_logic_bridge_dataFork_ready = 1'b1;
    end
  end

  assign LsuCachelessAxi4Plugin_logic_bridge_dataStage_payload_write = LsuCachelessAxi4Plugin_logic_bridge_dataFork_payload_write;
  assign LsuCachelessAxi4Plugin_logic_bridge_dataStage_payload_address = LsuCachelessAxi4Plugin_logic_bridge_dataFork_payload_address;
  assign LsuCachelessAxi4Plugin_logic_bridge_dataStage_payload_data = LsuCachelessAxi4Plugin_logic_bridge_dataFork_payload_data;
  assign LsuCachelessAxi4Plugin_logic_bridge_dataStage_payload_size = LsuCachelessAxi4Plugin_logic_bridge_dataFork_payload_size;
  assign LsuCachelessAxi4Plugin_logic_bridge_dataStage_payload_mask = LsuCachelessAxi4Plugin_logic_bridge_dataFork_payload_mask;
  assign LsuCachelessAxi4Plugin_logic_bridge_dataStage_payload_io = LsuCachelessAxi4Plugin_logic_bridge_dataFork_payload_io;
  assign LsuCachelessAxi4Plugin_logic_bridge_dataStage_payload_fromHart = LsuCachelessAxi4Plugin_logic_bridge_dataFork_payload_fromHart;
  assign LsuCachelessAxi4Plugin_logic_bridge_dataStage_payload_uopId = LsuCachelessAxi4Plugin_logic_bridge_dataFork_payload_uopId;
  assign LsuCachelessAxi4Plugin_logic_bridge_down_w_valid = LsuCachelessAxi4Plugin_logic_bridge_dataStage_valid;
  assign LsuCachelessAxi4Plugin_logic_bridge_dataStage_ready = LsuCachelessAxi4Plugin_logic_bridge_down_w_ready;
  assign LsuCachelessAxi4Plugin_logic_bridge_down_w_payload_last = 1'b1;
  assign LsuCachelessAxi4Plugin_logic_bridge_down_w_payload_data = LsuCachelessAxi4Plugin_logic_bridge_dataStage_payload_data;
  assign LsuCachelessAxi4Plugin_logic_bridge_down_w_payload_strb = LsuCachelessAxi4Plugin_logic_bridge_dataStage_payload_mask;
  always @(*) begin
    LsuPlugin_logic_bus_rsp_valid = LsuCachelessAxi4Plugin_logic_bridge_down_b_valid;
    if(LsuCachelessAxi4Plugin_logic_bridge_down_r_valid) begin
      LsuPlugin_logic_bus_rsp_valid = LsuCachelessAxi4Plugin_logic_bridge_down_r_valid;
    end
  end

  always @(*) begin
    LsuPlugin_logic_bus_rsp_payload_error = (! (LsuCachelessAxi4Plugin_logic_bridge_down_b_payload_resp == 2'b00));
    if(LsuCachelessAxi4Plugin_logic_bridge_down_r_valid) begin
      LsuPlugin_logic_bus_rsp_payload_error = (! (LsuCachelessAxi4Plugin_logic_bridge_down_r_payload_resp == 2'b00));
    end
  end

  assign LsuPlugin_logic_bus_rsp_payload_data = LsuCachelessAxi4Plugin_logic_bridge_down_r_payload_data;
  assign LsuCachelessAxi4Plugin_logic_bridge_down_r_ready = 1'b1;
  always @(*) begin
    LsuCachelessAxi4Plugin_logic_bridge_down_b_ready = 1'b1;
    if(LsuCachelessAxi4Plugin_logic_bridge_down_r_valid) begin
      LsuCachelessAxi4Plugin_logic_bridge_down_b_ready = 1'b0;
    end
  end

  assign LsuCachelessAxi4Plugin_logic_axi_ar_payload_addr = LsuCachelessAxi4Plugin_logic_bridge_down_arw_payload_addr;
  assign LsuCachelessAxi4Plugin_logic_axi_ar_payload_size = LsuCachelessAxi4Plugin_logic_bridge_down_arw_payload_size;
  assign LsuCachelessAxi4Plugin_logic_axi_ar_payload_cache = LsuCachelessAxi4Plugin_logic_bridge_down_arw_payload_cache;
  assign LsuCachelessAxi4Plugin_logic_axi_ar_payload_prot = LsuCachelessAxi4Plugin_logic_bridge_down_arw_payload_prot;
  assign LsuCachelessAxi4Plugin_logic_axi_aw_payload_addr = LsuCachelessAxi4Plugin_logic_bridge_down_arw_payload_addr;
  assign LsuCachelessAxi4Plugin_logic_axi_aw_payload_size = LsuCachelessAxi4Plugin_logic_bridge_down_arw_payload_size;
  assign LsuCachelessAxi4Plugin_logic_axi_aw_payload_cache = LsuCachelessAxi4Plugin_logic_bridge_down_arw_payload_cache;
  assign LsuCachelessAxi4Plugin_logic_axi_aw_payload_prot = LsuCachelessAxi4Plugin_logic_bridge_down_arw_payload_prot;
  assign LsuCachelessAxi4Plugin_logic_axi_ar_valid = (LsuCachelessAxi4Plugin_logic_bridge_down_arw_valid && (! LsuCachelessAxi4Plugin_logic_bridge_down_arw_payload_write));
  assign LsuCachelessAxi4Plugin_logic_axi_aw_valid = (LsuCachelessAxi4Plugin_logic_bridge_down_arw_valid && LsuCachelessAxi4Plugin_logic_bridge_down_arw_payload_write);
  assign LsuCachelessAxi4Plugin_logic_bridge_down_arw_ready = (LsuCachelessAxi4Plugin_logic_bridge_down_arw_payload_write ? LsuCachelessAxi4Plugin_logic_axi_aw_ready : LsuCachelessAxi4Plugin_logic_axi_ar_ready);
  assign LsuCachelessAxi4Plugin_logic_axi_w_valid = LsuCachelessAxi4Plugin_logic_bridge_down_w_valid;
  assign LsuCachelessAxi4Plugin_logic_bridge_down_w_ready = LsuCachelessAxi4Plugin_logic_axi_w_ready;
  assign LsuCachelessAxi4Plugin_logic_axi_w_payload_data = LsuCachelessAxi4Plugin_logic_bridge_down_w_payload_data;
  assign LsuCachelessAxi4Plugin_logic_axi_w_payload_strb = LsuCachelessAxi4Plugin_logic_bridge_down_w_payload_strb;
  assign LsuCachelessAxi4Plugin_logic_axi_w_payload_last = LsuCachelessAxi4Plugin_logic_bridge_down_w_payload_last;
  assign LsuCachelessAxi4Plugin_logic_bridge_down_r_valid = LsuCachelessAxi4Plugin_logic_axi_r_valid;
  assign LsuCachelessAxi4Plugin_logic_axi_r_ready = LsuCachelessAxi4Plugin_logic_bridge_down_r_ready;
  assign LsuCachelessAxi4Plugin_logic_bridge_down_r_payload_data = LsuCachelessAxi4Plugin_logic_axi_r_payload_data;
  assign LsuCachelessAxi4Plugin_logic_bridge_down_r_payload_resp = LsuCachelessAxi4Plugin_logic_axi_r_payload_resp;
  assign LsuCachelessAxi4Plugin_logic_bridge_down_r_payload_last = LsuCachelessAxi4Plugin_logic_axi_r_payload_last;
  assign LsuCachelessAxi4Plugin_logic_bridge_down_b_valid = LsuCachelessAxi4Plugin_logic_axi_b_valid;
  assign LsuCachelessAxi4Plugin_logic_axi_b_ready = LsuCachelessAxi4Plugin_logic_bridge_down_b_ready;
  assign LsuCachelessAxi4Plugin_logic_bridge_down_b_payload_resp = LsuCachelessAxi4Plugin_logic_axi_b_payload_resp;
  assign LsuPlugin_pmaBuilder_l1_addressBits = LsuPlugin_logic_onPma_cached_cmd_address;
  assign LsuPlugin_pmaBuilder_l1_argsBits = LsuPlugin_logic_onPma_cached_cmd_op;
  assign _zz_LsuPlugin_logic_onPma_cached_rsp_io = ((LsuPlugin_pmaBuilder_l1_addressBits & 32'h0) == 32'h0);
  assign LsuPlugin_pmaBuilder_l1_onTransfers_0_addressHit = _zz_LsuPlugin_pmaBuilder_l1_onTransfers_0_addressHit[0];
  assign LsuPlugin_pmaBuilder_l1_onTransfers_0_argsHit = (|((LsuPlugin_pmaBuilder_l1_argsBits & 1'b0) == 1'b0));
  assign LsuPlugin_pmaBuilder_l1_onTransfers_0_hit = (LsuPlugin_pmaBuilder_l1_onTransfers_0_argsHit && LsuPlugin_pmaBuilder_l1_onTransfers_0_addressHit);
  assign LsuPlugin_logic_onPma_cached_rsp_fault = (! ((|{((LsuPlugin_pmaBuilder_l1_addressBits & 32'hf8000000) == 32'h80000000),((LsuPlugin_pmaBuilder_l1_addressBits & 32'hf1000000) == 32'h0)}) && (|LsuPlugin_pmaBuilder_l1_onTransfers_0_hit)));
  assign LsuPlugin_logic_onPma_cached_rsp_io = (! _zz_LsuPlugin_logic_onPma_cached_rsp_io_1[0]);
  assign LsuPlugin_pmaBuilder_io_addressBits = LsuPlugin_logic_onPma_io_cmd_address;
  assign LsuPlugin_pmaBuilder_io_argsBits = {LsuPlugin_logic_onPma_io_cmd_size,LsuPlugin_logic_onPma_io_cmd_op};
  assign LsuPlugin_pmaBuilder_io_onTransfers_0_addressHit = _zz_LsuPlugin_pmaBuilder_io_onTransfers_0_addressHit[0];
  assign LsuPlugin_pmaBuilder_io_onTransfers_0_argsHit = (|((LsuPlugin_pmaBuilder_io_argsBits & 3'b000) == 3'b000));
  assign LsuPlugin_pmaBuilder_io_onTransfers_0_hit = (LsuPlugin_pmaBuilder_io_onTransfers_0_argsHit && LsuPlugin_pmaBuilder_io_onTransfers_0_addressHit);
  assign LsuPlugin_logic_onPma_io_rsp_fault = (! ((|{((LsuPlugin_pmaBuilder_io_addressBits & 32'he0000000) == 32'h40000000),{((LsuPlugin_pmaBuilder_io_addressBits & 32'he0000000) == 32'h20000000),{((LsuPlugin_pmaBuilder_io_addressBits & _zz_LsuPlugin_logic_onPma_io_rsp_fault) == 32'h60000000),{(_zz_LsuPlugin_logic_onPma_io_rsp_fault_1 == _zz_LsuPlugin_logic_onPma_io_rsp_fault_2),{_zz_LsuPlugin_logic_onPma_io_rsp_fault_3,{_zz_LsuPlugin_logic_onPma_io_rsp_fault_4,_zz_LsuPlugin_logic_onPma_io_rsp_fault_5}}}}}}) && (|LsuPlugin_pmaBuilder_io_onTransfers_0_hit)));
  assign LsuPlugin_logic_onPma_io_rsp_io = (! _zz_LsuPlugin_logic_onPma_io_rsp_io[0]);
  assign execute_ctrl2_down_early0_BranchPlugin_logic_alu_EQ_lane0 = ($signed(execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0) == $signed(execute_ctrl2_down_early0_SrcPlugin_SRC2_lane0));
  assign execute_ctrl2_down_early0_BranchPlugin_logic_alu_btb_BAD_TARGET_lane0 = (execute_ctrl2_down_Prediction_ALIGNED_JUMPED_PC_lane0 != execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0);
  assign early0_BranchPlugin_logic_alu_expectedMsb = (MmuPlugin_api_fetchTranslationEnable ? _zz_early0_BranchPlugin_logic_alu_expectedMsb[38] : 1'b0);
  assign _zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0 = _zz__zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0;
  assign execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0 = ((execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0 == BranchPlugin_BranchCtrlEnum_JALR) && (|{(_zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0[24] != early0_BranchPlugin_logic_alu_expectedMsb),{(_zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0[23] != early0_BranchPlugin_logic_alu_expectedMsb),{(_zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0[22] != early0_BranchPlugin_logic_alu_expectedMsb),{(_zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0_1 != early0_BranchPlugin_logic_alu_expectedMsb),{_zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0_2,{_zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0_3,_zz_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0_4}}}}}}));
  assign switch_Misc_l245_1 = execute_ctrl2_down_Decode_UOP_lane0[14 : 12];
  always @(*) begin
    casez(switch_Misc_l245_1)
      3'b000 : begin
        _zz_execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0 = execute_ctrl2_down_early0_BranchPlugin_logic_alu_EQ_lane0;
      end
      3'b001 : begin
        _zz_execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0 = (! execute_ctrl2_down_early0_BranchPlugin_logic_alu_EQ_lane0);
      end
      3'b1?1 : begin
        _zz_execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0 = (! execute_ctrl2_down_early0_SrcPlugin_LESS_lane0);
      end
      default : begin
        _zz_execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0 = execute_ctrl2_down_early0_SrcPlugin_LESS_lane0;
      end
    endcase
  end

  always @(*) begin
    case(execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0)
      BranchPlugin_BranchCtrlEnum_JALR : begin
        _zz_execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0_1 = 1'b1;
      end
      BranchPlugin_BranchCtrlEnum_JAL : begin
        _zz_execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0_1 = 1'b1;
      end
      default : begin
        _zz_execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0_1 = _zz_execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0;
      end
    endcase
  end

  assign execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0 = _zz_execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0_1;
  assign execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_btb_REAL_TARGET_lane0 = (execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0 ? execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0 : execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0);
  assign early0_BranchPlugin_logic_jumpLogic_wrongCond = (execute_ctrl2_down_Prediction_ALIGNED_JUMPED_lane0 != execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0);
  assign early0_BranchPlugin_logic_jumpLogic_needFix = ((early0_BranchPlugin_logic_jumpLogic_wrongCond || (execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0 && execute_ctrl2_down_early0_BranchPlugin_logic_alu_btb_BAD_TARGET_lane0)) || execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0);
  assign early0_BranchPlugin_logic_jumpLogic_doIt = ((execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_down_early0_BranchPlugin_SEL_lane0) && early0_BranchPlugin_logic_jumpLogic_needFix);
  assign early0_BranchPlugin_logic_jumpLogic_history_slice = execute_ctrl2_down_PC_lane0[1 : 1];
  assign early0_BranchPlugin_logic_jumpLogic_history_shifter = execute_ctrl2_down_Prediction_BRANCH_HISTORY_lane0;
  assign when_BranchPlugin_l213 = ((early0_BranchPlugin_logic_jumpLogic_history_slice < 1'b0) && execute_ctrl2_down_Prediction_ALIGNED_SLICES_BRANCH_lane0[0]);
  assign when_BranchPlugin_l218 = (execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0 == BranchPlugin_BranchCtrlEnum_B);
  assign early0_BranchPlugin_logic_jumpLogic_history_next = early0_BranchPlugin_logic_jumpLogic_history_shifter_2;
  assign early0_BranchPlugin_logic_jumpLogic_history_fetched = execute_ctrl2_down_Prediction_BRANCH_HISTORY_lane0;
  assign early0_BranchPlugin_logic_pcPort_valid = early0_BranchPlugin_logic_jumpLogic_doIt;
  assign early0_BranchPlugin_logic_pcPort_payload_fault = execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0;
  assign early0_BranchPlugin_logic_pcPort_payload_pc = execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_btb_REAL_TARGET_lane0;
  assign early0_BranchPlugin_logic_historyPort_valid = early0_BranchPlugin_logic_jumpLogic_doIt;
  assign early0_BranchPlugin_logic_historyPort_payload_history = early0_BranchPlugin_logic_jumpLogic_history_next;
  assign early0_BranchPlugin_logic_flushPort_valid = early0_BranchPlugin_logic_jumpLogic_doIt;
  assign early0_BranchPlugin_logic_flushPort_payload_uopId = execute_ctrl2_down_Decode_UOP_ID_lane0;
  assign early0_BranchPlugin_logic_flushPort_payload_self = 1'b0;
  assign execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_MISSALIGNED_lane0 = ((execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0[0 : 0] != 1'b0) && execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0);
  assign execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_IS_JAL_lane0 = (execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0 == BranchPlugin_BranchCtrlEnum_JAL);
  assign execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_IS_JALR_lane0 = (execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0 == BranchPlugin_BranchCtrlEnum_JALR);
  assign early0_BranchPlugin_logic_jumpLogic_rdLink = (|{(execute_ctrl2_down_Decode_UOP_lane0[11 : 7] == 5'h05),(execute_ctrl2_down_Decode_UOP_lane0[11 : 7] == 5'h01)});
  assign early0_BranchPlugin_logic_jumpLogic_rs1Link = (|{(execute_ctrl2_down_Decode_UOP_lane0[19 : 15] == 5'h05),(execute_ctrl2_down_Decode_UOP_lane0[19 : 15] == 5'h01)});
  assign early0_BranchPlugin_logic_jumpLogic_rdEquRs1 = (execute_ctrl2_down_Decode_UOP_lane0[11 : 7] == execute_ctrl2_down_Decode_UOP_lane0[19 : 15]);
  assign early0_BranchPlugin_logic_jumpLogic_learn_valid = (((execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_down_isReady) && (! execute_lane0_ctrls_2_upIsCancel)) && (|execute_ctrl2_down_early0_BranchPlugin_SEL_lane0));
  assign early0_BranchPlugin_logic_jumpLogic_learn_payload_taken = execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0;
  assign early0_BranchPlugin_logic_jumpLogic_learn_payload_pcTarget = execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0;
  assign early0_BranchPlugin_logic_jumpLogic_learn_payload_pcOnLastSlice = execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0;
  assign early0_BranchPlugin_logic_jumpLogic_learn_payload_isBranch = (execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0 == BranchPlugin_BranchCtrlEnum_B);
  assign early0_BranchPlugin_logic_jumpLogic_learn_payload_isPush = ((execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_IS_JAL_lane0 || execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_IS_JALR_lane0) && early0_BranchPlugin_logic_jumpLogic_rdLink);
  assign early0_BranchPlugin_logic_jumpLogic_learn_payload_isPop = (execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_IS_JALR_lane0 && (((! early0_BranchPlugin_logic_jumpLogic_rdLink) && early0_BranchPlugin_logic_jumpLogic_rs1Link) || ((early0_BranchPlugin_logic_jumpLogic_rdLink && early0_BranchPlugin_logic_jumpLogic_rs1Link) && (! early0_BranchPlugin_logic_jumpLogic_rdEquRs1))));
  assign early0_BranchPlugin_logic_jumpLogic_learn_payload_wasWrong = early0_BranchPlugin_logic_jumpLogic_needFix;
  assign early0_BranchPlugin_logic_jumpLogic_learn_payload_badPredictedTarget = execute_ctrl2_down_early0_BranchPlugin_logic_alu_btb_BAD_TARGET_lane0;
  assign early0_BranchPlugin_logic_jumpLogic_learn_payload_history = early0_BranchPlugin_logic_jumpLogic_history_fetched;
  assign early0_BranchPlugin_logic_jumpLogic_learn_payload_uopId = execute_ctrl2_down_Decode_UOP_ID_lane0;
  assign early0_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 = execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane0_0;
  assign early0_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_1 = execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane0_1;
  assign early0_BranchPlugin_logic_events_branchMiss = ((early0_BranchPlugin_logic_jumpLogic_learn_valid && early0_BranchPlugin_logic_jumpLogic_learn_payload_isBranch) && early0_BranchPlugin_logic_jumpLogic_learn_payload_wasWrong);
  assign early0_BranchPlugin_logic_events_branchCount = (early0_BranchPlugin_logic_jumpLogic_learn_valid && early0_BranchPlugin_logic_jumpLogic_learn_payload_isBranch);
  assign early0_BranchPlugin_logic_wb_valid = execute_ctrl2_down_early0_BranchPlugin_SEL_lane0;
  assign early0_BranchPlugin_logic_wb_payload = _zz_early0_BranchPlugin_logic_wb_payload;
  assign execute_ctrl2_COMPLETED_lane0_bypass = (execute_ctrl2_up_COMPLETED_lane0 || execute_ctrl2_down_COMPLETION_AT_2_lane0);
  assign execute_ctrl4_COMPLETED_lane0_bypass = (execute_ctrl4_up_COMPLETED_lane0 || execute_ctrl4_down_COMPLETION_AT_4_lane0);
  assign execute_ctrl3_COMPLETED_lane0_bypass = (execute_ctrl3_up_COMPLETED_lane0 || execute_ctrl3_down_COMPLETION_AT_3_lane0);
  assign execute_lane0_api_hartsInflight[0] = (|{(execute_ctrl4_up_LANE_SEL_lane0 && 1'b1),{(execute_ctrl3_up_LANE_SEL_lane0 && 1'b1),{(execute_ctrl2_up_LANE_SEL_lane0 && 1'b1),(execute_ctrl1_up_LANE_SEL_lane0 && 1'b1)}}});
  assign LearnPlugin_logic_buffered_0_valid = early0_BranchPlugin_logic_jumpLogic_learn_valid;
  assign early0_BranchPlugin_logic_jumpLogic_learn_ready = LearnPlugin_logic_buffered_0_ready;
  assign LearnPlugin_logic_buffered_0_payload_pcOnLastSlice = early0_BranchPlugin_logic_jumpLogic_learn_payload_pcOnLastSlice;
  assign LearnPlugin_logic_buffered_0_payload_pcTarget = early0_BranchPlugin_logic_jumpLogic_learn_payload_pcTarget;
  assign LearnPlugin_logic_buffered_0_payload_taken = early0_BranchPlugin_logic_jumpLogic_learn_payload_taken;
  assign LearnPlugin_logic_buffered_0_payload_isBranch = early0_BranchPlugin_logic_jumpLogic_learn_payload_isBranch;
  assign LearnPlugin_logic_buffered_0_payload_isPush = early0_BranchPlugin_logic_jumpLogic_learn_payload_isPush;
  assign LearnPlugin_logic_buffered_0_payload_isPop = early0_BranchPlugin_logic_jumpLogic_learn_payload_isPop;
  assign LearnPlugin_logic_buffered_0_payload_wasWrong = early0_BranchPlugin_logic_jumpLogic_learn_payload_wasWrong;
  assign LearnPlugin_logic_buffered_0_payload_badPredictedTarget = early0_BranchPlugin_logic_jumpLogic_learn_payload_badPredictedTarget;
  assign LearnPlugin_logic_buffered_0_payload_history = early0_BranchPlugin_logic_jumpLogic_learn_payload_history;
  assign LearnPlugin_logic_buffered_0_payload_uopId = early0_BranchPlugin_logic_jumpLogic_learn_payload_uopId;
  assign LearnPlugin_logic_buffered_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 = early0_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  assign LearnPlugin_logic_buffered_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_1 = early0_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  assign LearnPlugin_logic_buffered_0_ready = streamArbiter_5_io_inputs_0_ready;
  assign LearnPlugin_logic_arbitrated_valid = streamArbiter_5_io_output_valid;
  assign LearnPlugin_logic_arbitrated_payload_pcOnLastSlice = streamArbiter_5_io_output_payload_pcOnLastSlice;
  assign LearnPlugin_logic_arbitrated_payload_pcTarget = streamArbiter_5_io_output_payload_pcTarget;
  assign LearnPlugin_logic_arbitrated_payload_taken = streamArbiter_5_io_output_payload_taken;
  assign LearnPlugin_logic_arbitrated_payload_isBranch = streamArbiter_5_io_output_payload_isBranch;
  assign LearnPlugin_logic_arbitrated_payload_isPush = streamArbiter_5_io_output_payload_isPush;
  assign LearnPlugin_logic_arbitrated_payload_isPop = streamArbiter_5_io_output_payload_isPop;
  assign LearnPlugin_logic_arbitrated_payload_wasWrong = streamArbiter_5_io_output_payload_wasWrong;
  assign LearnPlugin_logic_arbitrated_payload_badPredictedTarget = streamArbiter_5_io_output_payload_badPredictedTarget;
  assign LearnPlugin_logic_arbitrated_payload_history = streamArbiter_5_io_output_payload_history;
  assign LearnPlugin_logic_arbitrated_payload_uopId = streamArbiter_5_io_output_payload_uopId;
  assign LearnPlugin_logic_arbitrated_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 = streamArbiter_5_io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  assign LearnPlugin_logic_arbitrated_payload_ctx_GSharePlugin_GSHARE_COUNTER_1 = streamArbiter_5_io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  assign LearnPlugin_logic_arbitrated_ready = 1'b1;
  assign LearnPlugin_logic_arbitrated_toFlow_valid = LearnPlugin_logic_arbitrated_valid;
  assign LearnPlugin_logic_arbitrated_toFlow_payload_pcOnLastSlice = LearnPlugin_logic_arbitrated_payload_pcOnLastSlice;
  assign LearnPlugin_logic_arbitrated_toFlow_payload_pcTarget = LearnPlugin_logic_arbitrated_payload_pcTarget;
  assign LearnPlugin_logic_arbitrated_toFlow_payload_taken = LearnPlugin_logic_arbitrated_payload_taken;
  assign LearnPlugin_logic_arbitrated_toFlow_payload_isBranch = LearnPlugin_logic_arbitrated_payload_isBranch;
  assign LearnPlugin_logic_arbitrated_toFlow_payload_isPush = LearnPlugin_logic_arbitrated_payload_isPush;
  assign LearnPlugin_logic_arbitrated_toFlow_payload_isPop = LearnPlugin_logic_arbitrated_payload_isPop;
  assign LearnPlugin_logic_arbitrated_toFlow_payload_wasWrong = LearnPlugin_logic_arbitrated_payload_wasWrong;
  assign LearnPlugin_logic_arbitrated_toFlow_payload_badPredictedTarget = LearnPlugin_logic_arbitrated_payload_badPredictedTarget;
  assign LearnPlugin_logic_arbitrated_toFlow_payload_history = LearnPlugin_logic_arbitrated_payload_history;
  assign LearnPlugin_logic_arbitrated_toFlow_payload_uopId = LearnPlugin_logic_arbitrated_payload_uopId;
  assign LearnPlugin_logic_arbitrated_toFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 = LearnPlugin_logic_arbitrated_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  assign LearnPlugin_logic_arbitrated_toFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_1 = LearnPlugin_logic_arbitrated_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  assign LearnPlugin_logic_learn_valid = LearnPlugin_logic_arbitrated_toFlow_valid;
  assign LearnPlugin_logic_learn_payload_pcOnLastSlice = LearnPlugin_logic_arbitrated_toFlow_payload_pcOnLastSlice;
  assign LearnPlugin_logic_learn_payload_pcTarget = LearnPlugin_logic_arbitrated_toFlow_payload_pcTarget;
  assign LearnPlugin_logic_learn_payload_taken = LearnPlugin_logic_arbitrated_toFlow_payload_taken;
  assign LearnPlugin_logic_learn_payload_isBranch = LearnPlugin_logic_arbitrated_toFlow_payload_isBranch;
  assign LearnPlugin_logic_learn_payload_isPush = LearnPlugin_logic_arbitrated_toFlow_payload_isPush;
  assign LearnPlugin_logic_learn_payload_isPop = LearnPlugin_logic_arbitrated_toFlow_payload_isPop;
  assign LearnPlugin_logic_learn_payload_wasWrong = LearnPlugin_logic_arbitrated_toFlow_payload_wasWrong;
  assign LearnPlugin_logic_learn_payload_badPredictedTarget = LearnPlugin_logic_arbitrated_toFlow_payload_badPredictedTarget;
  assign LearnPlugin_logic_learn_payload_history = LearnPlugin_logic_arbitrated_toFlow_payload_history;
  assign LearnPlugin_logic_learn_payload_uopId = LearnPlugin_logic_arbitrated_toFlow_payload_uopId;
  assign LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 = LearnPlugin_logic_arbitrated_toFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  assign LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_1 = LearnPlugin_logic_arbitrated_toFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  assign when_DecoderPlugin_l143 = (decode_ctrls_1_up_isMoving && 1'b1);
  assign DecoderPlugin_logic_interrupt_async = PrivilegedPlugin_logic_harts_0_int_pending;
  assign when_DecoderPlugin_l151 = (((! decode_ctrls_1_up_valid) || decode_ctrls_1_up_ready) || decode_ctrls_1_up_isCanceling);
  assign decode_ctrls_1_down_RS1_ENABLE_0 = _zz_decode_ctrls_1_down_RS1_ENABLE_0[0];
  assign decode_ctrls_1_down_RS1_PHYS_0 = _zz_decode_ctrls_1_down_RS1_PHYS_0[4 : 0];
  assign decode_ctrls_1_down_RS2_ENABLE_0 = _zz_decode_ctrls_1_down_RS2_ENABLE_0[0];
  assign decode_ctrls_1_down_RS2_PHYS_0 = _zz_decode_ctrls_1_down_RS2_PHYS_0[4 : 0];
  always @(*) begin
    decode_ctrls_1_down_RD_ENABLE_0 = _zz_decode_ctrls_1_down_RD_ENABLE_0[0];
    if(when_DecoderPlugin_l247) begin
      decode_ctrls_1_down_RD_ENABLE_0 = 1'b0;
    end
  end

  assign decode_ctrls_1_down_RD_PHYS_0 = _zz_decode_ctrls_1_down_RD_PHYS_0[4 : 0];
  always @(*) begin
    decode_ctrls_1_down_Decode_LEGAL_0 = ((|{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000005f) == 32'h00000017),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000007f) == 32'h0000006f),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & _zz_decode_ctrls_1_down_Decode_LEGAL_0) == 32'h00000003),{(_zz_decode_ctrls_1_down_Decode_LEGAL_0_1 == _zz_decode_ctrls_1_down_Decode_LEGAL_0_2),{_zz_decode_ctrls_1_down_Decode_LEGAL_0_3,{_zz_decode_ctrls_1_down_Decode_LEGAL_0_4,_zz_decode_ctrls_1_down_Decode_LEGAL_0_5}}}}}}) && (! decode_ctrls_1_down_Decode_DECOMPRESSION_FAULT_0));
    if(when_DecoderPlugin_l187) begin
      decode_ctrls_1_down_Decode_LEGAL_0 = 1'b0;
    end
    if(when_DecoderPlugin_l187_1) begin
      decode_ctrls_1_down_Decode_LEGAL_0 = 1'b0;
    end
  end

  assign when_DecoderPlugin_l187 = (LsuPlugin_logic_cbmCsr_menvcfg_privLower && ((decode_ctrls_1_down_AguPlugin_INVALIDATE_0 && (LsuPlugin_logic_cbmCsr_menvcfg_cbie == 2'b00)) || ((decode_ctrls_1_down_AguPlugin_CLEAN_0 && (LsuPlugin_logic_cbmCsr_menvcfg_cbcfe == 1'b0)) && LsuPlugin_logic_cbmCsr_menvcfg_privLower)));
  assign when_DecoderPlugin_l187_1 = (LsuPlugin_logic_cbmCsr_senvcfg_privLower && ((decode_ctrls_1_down_AguPlugin_INVALIDATE_0 && (LsuPlugin_logic_cbmCsr_senvcfg_cbie == 2'b00)) || ((decode_ctrls_1_down_AguPlugin_CLEAN_0 && (LsuPlugin_logic_cbmCsr_senvcfg_cbcfe == 1'b0)) && LsuPlugin_logic_cbmCsr_senvcfg_privLower)));
  assign DecoderPlugin_logic_laneLogic_0_interruptPending = DecoderPlugin_logic_interrupt_buffered[0];
  always @(*) begin
    DecoderPlugin_logic_laneLogic_0_trapPort_valid = 1'b0;
    if(when_DecoderPlugin_l229) begin
      DecoderPlugin_logic_laneLogic_0_trapPort_valid = ((! decode_ctrls_1_up_TRAP_0) || DecoderPlugin_logic_laneLogic_0_interruptPending);
      if(DecoderPlugin_logic_laneLogic_0_fixer_doIt) begin
        DecoderPlugin_logic_laneLogic_0_trapPort_valid = 1'b1;
      end
    end
  end

  always @(*) begin
    DecoderPlugin_logic_laneLogic_0_trapPort_payload_exception = 1'b1;
    if(DecoderPlugin_logic_laneLogic_0_fixer_doIt) begin
      DecoderPlugin_logic_laneLogic_0_trapPort_payload_exception = 1'b0;
    end
    if(DecoderPlugin_logic_laneLogic_0_interruptPending) begin
      DecoderPlugin_logic_laneLogic_0_trapPort_payload_exception = 1'b0;
    end
  end

  assign DecoderPlugin_logic_laneLogic_0_trapPort_payload_tval = {7'd0, decode_ctrls_1_down_Decode_INSTRUCTION_RAW_0};
  always @(*) begin
    DecoderPlugin_logic_laneLogic_0_trapPort_payload_code = 4'b0010;
    if(DecoderPlugin_logic_laneLogic_0_fixer_doIt) begin
      DecoderPlugin_logic_laneLogic_0_trapPort_payload_code = 4'b0100;
    end
    if(DecoderPlugin_logic_laneLogic_0_interruptPending) begin
      DecoderPlugin_logic_laneLogic_0_trapPort_payload_code = 4'b0000;
    end
  end

  assign DecoderPlugin_logic_laneLogic_0_trapPort_payload_laneAge = 1'b0;
  assign DecoderPlugin_logic_laneLogic_0_trapPort_payload_arg = 3'b000;
  assign DecoderPlugin_logic_laneLogic_0_fixer_isJb = _zz_DecoderPlugin_logic_laneLogic_0_fixer_isJb[0];
  assign DecoderPlugin_logic_laneLogic_0_fixer_doIt = (decode_ctrls_1_up_LANE_SEL_0 && ((decode_ctrls_1_down_Prediction_ALIGNED_JUMPED_0 && (! DecoderPlugin_logic_laneLogic_0_fixer_isJb)) || decode_ctrls_1_down_Prediction_ALIGN_REDO_0));
  assign when_CtrlLaneApi_l50_1 = (decode_ctrls_1_up_isReady || decode_ctrls_1_lane0_upIsCancel);
  assign DecoderPlugin_logic_laneLogic_0_completionPort_valid = ((decode_ctrls_1_up_LANE_SEL_0 && decode_ctrls_1_down_TRAP_0) && (decode_ctrls_1_up_LANE_SEL_0 && (! decode_ctrls_1_up_LANE_SEL_0_regNext)));
  assign DecoderPlugin_logic_laneLogic_0_completionPort_payload_uopId = decode_ctrls_1_down_Decode_UOP_ID_0;
  assign DecoderPlugin_logic_laneLogic_0_completionPort_payload_trap = 1'b1;
  assign DecoderPlugin_logic_laneLogic_0_completionPort_payload_commit = 1'b0;
  assign when_DecoderPlugin_l229 = (decode_ctrls_1_up_LANE_SEL_0 && (((! decode_ctrls_1_down_Decode_LEGAL_0) || DecoderPlugin_logic_laneLogic_0_interruptPending) || DecoderPlugin_logic_laneLogic_0_fixer_doIt));
  assign DecoderPlugin_logic_laneLogic_0_flushPort_valid = (decode_ctrls_1_up_LANE_SEL_0 && decode_ctrls_1_down_TRAP_0);
  assign DecoderPlugin_logic_laneLogic_0_flushPort_payload_uopId = decode_ctrls_1_down_Decode_UOP_ID_0;
  assign DecoderPlugin_logic_laneLogic_0_flushPort_payload_self = 1'b0;
  assign when_DecoderPlugin_l247 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0[11 : 7] == 5'h0) && (|1'b1));
  assign decode_ctrls_1_down_Decode_UOP_0 = decode_ctrls_1_down_Decode_INSTRUCTION_0;
  assign DecoderPlugin_logic_laneLogic_0_uopIdBase = DecoderPlugin_logic_harts_0_uopId;
  assign decode_ctrls_1_down_Decode_UOP_ID_0 = (DecoderPlugin_logic_laneLogic_0_uopIdBase + 16'h0);
  assign DispatchPlugin_logic_trapPendings[0] = 1'b0;
  assign DispatchPlugin_logic_candidates_0_moving = (((! DispatchPlugin_logic_candidates_0_ctx_valid) || DispatchPlugin_logic_candidates_0_fire) || DispatchPlugin_logic_candidates_0_cancel);
  assign DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard = (DispatchPlugin_logic_candidates_0_ctx_hm_RS1_ENABLE && (|{((((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 && execute_ctrl2_up_RD_ENABLE_lane0) && (execute_ctrl2_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS1_PHYS)) && 1'b1) && (! execute_ctrl2_down_BYPASSED_AT_3_lane0)),((((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 && execute_ctrl1_up_RD_ENABLE_lane0) && (execute_ctrl1_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS1_PHYS)) && 1'b1) && (! execute_ctrl1_down_BYPASSED_AT_2_lane0))}));
  assign DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard = (DispatchPlugin_logic_candidates_0_ctx_hm_RS2_ENABLE && (|{((((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 && execute_ctrl2_up_RD_ENABLE_lane0) && (execute_ctrl2_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS2_PHYS)) && 1'b1) && (! execute_ctrl2_down_BYPASSED_AT_3_lane0)),((((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 && execute_ctrl1_up_RD_ENABLE_lane0) && (execute_ctrl1_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS2_PHYS)) && 1'b1) && (! execute_ctrl1_down_BYPASSED_AT_2_lane0))}));
  assign DispatchPlugin_logic_candidates_0_rsHazards[0] = (|{DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard,DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard});
  assign DispatchPlugin_logic_reservationChecker_0_onLl_0_hit = 1'b0;
  assign DispatchPlugin_logic_candidates_0_reservationHazards[0] = DispatchPlugin_logic_reservationChecker_0_onLl_0_hit;
  assign DispatchPlugin_logic_flushChecker_0_executeCheck_0_hits_0 = (|{(((DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_4 && execute_ctrl1_up_LANE_SEL_lane0) && 1'b1) && execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane0),(((DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_3 && execute_ctrl1_up_LANE_SEL_lane0) && 1'b1) && execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane0)});
  assign DispatchPlugin_logic_flushChecker_0_executeCheck_0_hits_1 = (|(((DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_3 && execute_ctrl2_up_LANE_SEL_lane0) && 1'b1) && execute_ctrl2_down_MAY_FLUSH_PRECISE_3_lane0));
  assign DispatchPlugin_logic_flushChecker_0_oldersHazard = 1'b0;
  assign DispatchPlugin_logic_candidates_0_flushHazards = ((|{DispatchPlugin_logic_flushChecker_0_executeCheck_0_hits_1,DispatchPlugin_logic_flushChecker_0_executeCheck_0_hits_0}) || (DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES && DispatchPlugin_logic_flushChecker_0_oldersHazard));
  assign DispatchPlugin_logic_fenceChecker_olderInflights = (|execute_lane0_api_hartsInflight[0]);
  assign DispatchPlugin_logic_candidates_0_fenceOlderHazards = (DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_FENCE_OLDER && (DispatchPlugin_logic_fenceChecker_olderInflights[0] || 1'b0));
  always @(*) begin
    decode_ctrls_1_down_ready = 1'b1;
    if(when_DispatchPlugin_l368) begin
      decode_ctrls_1_down_ready = 1'b0;
    end
  end

  assign DispatchPlugin_logic_feeds_0_sending = DispatchPlugin_logic_candidates_0_fire;
  assign DispatchPlugin_logic_candidates_0_cancel = decode_ctrls_1_lane0_upIsCancel;
  assign DispatchPlugin_logic_candidates_0_ctx_valid = ((decode_ctrls_1_up_isValid && decode_ctrls_1_up_LANE_SEL_0) && (! DispatchPlugin_logic_feeds_0_sent));
  always @(*) begin
    DispatchPlugin_logic_candidates_0_ctx_laneLayerHits = decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0;
    if(decode_ctrls_1_down_TRAP_0) begin
      DispatchPlugin_logic_candidates_0_ctx_laneLayerHits = 1'b1;
    end
  end

  assign DispatchPlugin_logic_candidates_0_ctx_uop = decode_ctrls_1_down_Decode_UOP_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_JUMPED = decode_ctrls_1_down_Prediction_ALIGNED_JUMPED_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_JUMPED_PC = decode_ctrls_1_down_Prediction_ALIGNED_JUMPED_PC_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_SLICES_TAKEN = decode_ctrls_1_down_Prediction_ALIGNED_SLICES_TAKEN_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_SLICES_BRANCH = decode_ctrls_1_down_Prediction_ALIGNED_SLICES_BRANCH_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_0 = decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_1 = decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0_1;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_BRANCH_HISTORY = decode_ctrls_1_down_Prediction_BRANCH_HISTORY_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_FENCE_OLDER = decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_MAY_FLUSH = decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_DONT_FLUSH = decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES = decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_Decode_INSTRUCTION_SLICE_COUNT = decode_ctrls_1_down_Decode_INSTRUCTION_SLICE_COUNT_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_3 = decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_4 = decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_PC = decode_ctrls_1_down_PC_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_TRAP = decode_ctrls_1_down_TRAP_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_Decode_UOP_ID = decode_ctrls_1_down_Decode_UOP_ID_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_RS1_ENABLE = decode_ctrls_1_down_RS1_ENABLE_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_RS1_PHYS = decode_ctrls_1_down_RS1_PHYS_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_RS2_ENABLE = decode_ctrls_1_down_RS2_ENABLE_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_RS2_PHYS = decode_ctrls_1_down_RS2_PHYS_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_RD_ENABLE = decode_ctrls_1_down_RD_ENABLE_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_RD_PHYS = decode_ctrls_1_down_RD_PHYS_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 = decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 = decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0;
  assign when_DispatchPlugin_l368 = ((decode_ctrls_1_up_LANE_SEL_0 && (! DispatchPlugin_logic_feeds_0_sent)) && (! DispatchPlugin_logic_candidates_0_fire));
  assign DispatchPlugin_logic_scheduler_eusFree_0 = 1'b1;
  assign DispatchPlugin_logic_scheduler_hartFree_0 = 1'b1;
  assign DispatchPlugin_logic_scheduler_arbiters_0_candHazard = 1'b0;
  assign DispatchPlugin_logic_scheduler_arbiters_0_layersHits = (((DispatchPlugin_logic_candidates_0_ctx_laneLayerHits & (~ DispatchPlugin_logic_candidates_0_rsHazards)) & (~ DispatchPlugin_logic_candidates_0_reservationHazards)) & DispatchPlugin_logic_scheduler_eusFree_0[0]);
  assign DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_0 = DispatchPlugin_logic_scheduler_arbiters_0_layersHits[0];
  assign _zz_DispatchPlugin_logic_scheduler_arbiters_0_layerOh[0] = (DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_0 && (! 1'b0));
  assign DispatchPlugin_logic_scheduler_arbiters_0_layerOh = _zz_DispatchPlugin_logic_scheduler_arbiters_0_layerOh;
  assign DispatchPlugin_logic_scheduler_arbiters_0_eusOh = (|DispatchPlugin_logic_scheduler_arbiters_0_layerOh[0]);
  assign DispatchPlugin_logic_scheduler_arbiters_0_doIt = (((((DispatchPlugin_logic_candidates_0_ctx_valid && (! DispatchPlugin_logic_candidates_0_flushHazards)) && (! DispatchPlugin_logic_candidates_0_fenceOlderHazards)) && (|DispatchPlugin_logic_scheduler_arbiters_0_layerOh)) && DispatchPlugin_logic_scheduler_hartFree_0[0]) && (! DispatchPlugin_logic_scheduler_arbiters_0_candHazard));
  assign DispatchPlugin_logic_scheduler_eusFree_1 = (DispatchPlugin_logic_scheduler_eusFree_0 & ((! DispatchPlugin_logic_scheduler_arbiters_0_doIt) ? 1'b1 : (~ DispatchPlugin_logic_scheduler_arbiters_0_eusOh)));
  assign DispatchPlugin_logic_scheduler_hartFree_1 = (DispatchPlugin_logic_scheduler_hartFree_0 & (((! DispatchPlugin_logic_candidates_0_ctx_valid) || DispatchPlugin_logic_scheduler_arbiters_0_doIt) ? 1'b1 : (~ 1'b1)));
  assign DispatchPlugin_logic_candidates_0_fire = ((DispatchPlugin_logic_scheduler_arbiters_0_doIt && (! execute_freeze_valid)) && (! DispatchPlugin_api_haltDispatch));
  assign DispatchPlugin_logic_inserter_0_oh = (DispatchPlugin_logic_scheduler_arbiters_0_doIt && DispatchPlugin_logic_scheduler_arbiters_0_eusOh[0]);
  assign DispatchPlugin_logic_inserter_0_trap = DispatchPlugin_logic_candidates_0_ctx_hm_TRAP;
  assign execute_ctrl0_up_LANE_SEL_lane0 = (((|DispatchPlugin_logic_inserter_0_oh) && (! DispatchPlugin_logic_candidates_0_cancel)) && (! DispatchPlugin_api_haltDispatch));
  assign execute_ctrl0_up_Decode_UOP_lane0 = DispatchPlugin_logic_candidates_0_ctx_uop;
  assign execute_ctrl0_up_Prediction_ALIGNED_JUMPED_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_JUMPED;
  assign execute_ctrl0_up_Prediction_ALIGNED_JUMPED_PC_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_JUMPED_PC;
  assign execute_ctrl0_up_Prediction_ALIGNED_SLICES_TAKEN_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_SLICES_TAKEN;
  assign execute_ctrl0_up_Prediction_ALIGNED_SLICES_BRANCH_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_SLICES_BRANCH;
  assign execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0 = DispatchPlugin_logic_candidates_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_0;
  assign execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_1 = DispatchPlugin_logic_candidates_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_1;
  assign execute_ctrl0_up_Prediction_BRANCH_HISTORY_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_BRANCH_HISTORY;
  assign execute_ctrl0_up_DispatchPlugin_FENCE_OLDER_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_FENCE_OLDER;
  always @(*) begin
    execute_ctrl0_up_DispatchPlugin_MAY_FLUSH_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_MAY_FLUSH;
    if(when_DispatchPlugin_l439) begin
      execute_ctrl0_up_DispatchPlugin_MAY_FLUSH_lane0 = 1'b0;
    end
  end

  assign execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_DONT_FLUSH;
  assign execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_FROM_LANES_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES;
  assign execute_ctrl0_up_Decode_INSTRUCTION_SLICE_COUNT_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_Decode_INSTRUCTION_SLICE_COUNT;
  assign execute_ctrl0_up_DONT_FLUSH_PRECISE_3_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_3;
  assign execute_ctrl0_up_DONT_FLUSH_PRECISE_4_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_4;
  assign execute_ctrl0_up_PC_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_PC;
  assign execute_ctrl0_up_TRAP_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_TRAP;
  assign execute_ctrl0_up_Decode_UOP_ID_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_Decode_UOP_ID;
  assign execute_ctrl0_up_RS1_ENABLE_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_RS1_ENABLE;
  assign execute_ctrl0_up_RS1_PHYS_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_RS1_PHYS;
  assign execute_ctrl0_up_RS2_ENABLE_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_RS2_ENABLE;
  assign execute_ctrl0_up_RS2_PHYS_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_RS2_PHYS;
  always @(*) begin
    execute_ctrl0_up_RD_ENABLE_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_RD_ENABLE;
    if(when_DispatchPlugin_l439) begin
      execute_ctrl0_up_RD_ENABLE_lane0 = 1'b0;
    end
  end

  assign execute_ctrl0_up_RD_PHYS_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_RD_PHYS;
  assign execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0;
  assign execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0;
  assign when_DispatchPlugin_l439 = ((! execute_ctrl0_up_LANE_SEL_lane0) || DispatchPlugin_logic_inserter_0_trap);
  assign execute_ctrl0_up_COMPLETED_lane0 = DispatchPlugin_logic_inserter_0_trap;
  assign DispatchPlugin_logic_inserter_0_layerOhUnfiltred = (DispatchPlugin_logic_inserter_0_oh[0] ? DispatchPlugin_logic_scheduler_arbiters_0_layerOh : 1'b0);
  assign DispatchPlugin_logic_inserter_0_layer_0_1 = DispatchPlugin_logic_inserter_0_layerOhUnfiltred[0];
  assign DispatchPlugin_logic_events_frontendStall = (DispatchPlugin_logic_candidates_0_ctx_valid == 1'b0);
  assign DispatchPlugin_logic_events_backendStall = ((|DispatchPlugin_logic_candidates_0_ctx_valid) && (DispatchPlugin_logic_candidates_0_fire == 1'b0));
  assign _zz_CsrRamPlugin_csrMapper_ramAddress = CsrAccessPlugin_bus_decode_address;
  assign CsrRamPlugin_csrMapper_ramAddress = {(|{(_zz_CsrRamPlugin_csrMapper_ramAddress_1 == _zz_CsrRamPlugin_csrMapper_ramAddress_2),(_zz_CsrRamPlugin_csrMapper_ramAddress_3 == _zz_CsrRamPlugin_csrMapper_ramAddress_4)}),{(|{_zz_CsrRamPlugin_csrMapper_ramAddress_5,{_zz_CsrRamPlugin_csrMapper_ramAddress_6,_zz_CsrRamPlugin_csrMapper_ramAddress_8}}),{(|_zz_CsrRamPlugin_csrMapper_ramAddress_10),(|{_zz_CsrRamPlugin_csrMapper_ramAddress_11,_zz_CsrRamPlugin_csrMapper_ramAddress_13})}}};
  always @(*) begin
    CsrRamPlugin_csrMapper_withRead = 1'b0;
    if(when_CsrAccessPlugin_l258) begin
      CsrRamPlugin_csrMapper_withRead = 1'b1;
    end
  end

  assign CsrRamPlugin_csrMapper_read_valid = (CsrRamPlugin_csrMapper_withRead && (! CsrRamPlugin_api_holdRead));
  assign CsrRamPlugin_csrMapper_read_address = CsrRamPlugin_csrMapper_ramAddress;
  assign when_CsrRamPlugin_l90 = (CsrRamPlugin_csrMapper_withRead && (! CsrRamPlugin_csrMapper_read_ready));
  always @(*) begin
    CsrRamPlugin_csrMapper_doWrite = 1'b0;
    if(when_CsrAccessPlugin_l349_2) begin
      CsrRamPlugin_csrMapper_doWrite = 1'b1;
    end
  end

  assign when_CsrRamPlugin_l97 = (CsrRamPlugin_csrMapper_write_valid && CsrRamPlugin_csrMapper_write_ready);
  assign CsrRamPlugin_csrMapper_write_valid = ((CsrRamPlugin_csrMapper_doWrite && (! CsrRamPlugin_csrMapper_fired)) && (! CsrRamPlugin_api_holdWrite));
  assign CsrRamPlugin_csrMapper_write_address = CsrRamPlugin_csrMapper_ramAddress;
  assign CsrRamPlugin_csrMapper_write_data = CsrAccessPlugin_bus_write_bits;
  assign when_CsrRamPlugin_l101 = ((CsrRamPlugin_csrMapper_doWrite && (! CsrRamPlugin_csrMapper_fired)) && (! CsrRamPlugin_csrMapper_write_ready));
  assign _zz_GSharePlugin_logic_onLearn_hash = LearnPlugin_logic_learn_payload_pcOnLastSlice[14 : 2];
  assign GSharePlugin_logic_onLearn_hash = ({_zz_GSharePlugin_logic_onLearn_hash[0],{_zz_GSharePlugin_logic_onLearn_hash[1],{_zz_GSharePlugin_logic_onLearn_hash[2],{_zz_GSharePlugin_logic_onLearn_hash[3],{_zz_GSharePlugin_logic_onLearn_hash[4],{_zz_GSharePlugin_logic_onLearn_hash[5],{_zz_GSharePlugin_logic_onLearn_hash_1,{_zz_GSharePlugin_logic_onLearn_hash_2,_zz_GSharePlugin_logic_onLearn_hash_3}}}}}}}} ^ _zz_GSharePlugin_logic_onLearn_hash_4);
  assign GSharePlugin_logic_onLearn_incrValue = (LearnPlugin_logic_learn_payload_taken ? 2'b01 : 2'b11);
  always @(*) begin
    GSharePlugin_logic_onLearn_overflow = 1'b0;
    if(when_GSharePlugin_l119) begin
      GSharePlugin_logic_onLearn_overflow = 1'b1;
    end
    if(when_GSharePlugin_l119_1) begin
      GSharePlugin_logic_onLearn_overflow = 1'b1;
    end
  end

  assign GSharePlugin_logic_onLearn_updated_0 = (LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 + ((LearnPlugin_logic_learn_payload_pcOnLastSlice[1 : 1] == 1'b0) ? GSharePlugin_logic_onLearn_incrValue : 2'b00));
  assign when_GSharePlugin_l119 = (((LearnPlugin_logic_learn_payload_taken && LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_0[1]) && (! GSharePlugin_logic_onLearn_updated_0[1])) || (((! LearnPlugin_logic_learn_payload_taken) && (! LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_0[1])) && GSharePlugin_logic_onLearn_updated_0[1]));
  assign GSharePlugin_logic_onLearn_updated_1 = (LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_1 + ((LearnPlugin_logic_learn_payload_pcOnLastSlice[1 : 1] == 1'b1) ? GSharePlugin_logic_onLearn_incrValue : 2'b00));
  assign when_GSharePlugin_l119_1 = (((LearnPlugin_logic_learn_payload_taken && LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_1[1]) && (! GSharePlugin_logic_onLearn_updated_1[1])) || (((! LearnPlugin_logic_learn_payload_taken) && (! LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_1[1])) && GSharePlugin_logic_onLearn_updated_1[1]));
  assign GSharePlugin_logic_mem_write_valid = ((LearnPlugin_logic_learn_valid && LearnPlugin_logic_learn_payload_isBranch) && (! GSharePlugin_logic_onLearn_overflow));
  assign GSharePlugin_logic_mem_write_payload_address = GSharePlugin_logic_onLearn_hash;
  assign GSharePlugin_logic_mem_write_payload_data_0 = GSharePlugin_logic_onLearn_updated_0;
  assign GSharePlugin_logic_mem_write_payload_data_1 = GSharePlugin_logic_onLearn_updated_1;
  assign BtbPlugin_logic_onLearn_hash = LearnPlugin_logic_learn_payload_pcOnLastSlice[26 : 11];
  always @(*) begin
    BtbPlugin_logic_memWrite_valid = (LearnPlugin_logic_learn_valid && (LearnPlugin_logic_learn_payload_badPredictedTarget && LearnPlugin_logic_learn_payload_taken));
    if(DecoderPlugin_logic_forgetPort_valid) begin
      BtbPlugin_logic_memWrite_valid = DecoderPlugin_logic_forgetPort_valid;
    end
  end

  always @(*) begin
    BtbPlugin_logic_memWrite_payload_address = _zz_BtbPlugin_logic_memWrite_payload_address[8:0];
    if(DecoderPlugin_logic_forgetPort_valid) begin
      BtbPlugin_logic_memWrite_payload_address = _zz_BtbPlugin_logic_memWrite_payload_address_1[8:0];
    end
  end

  always @(*) begin
    BtbPlugin_logic_memWrite_payload_mask = 1'b1;
    if(DecoderPlugin_logic_forgetPort_valid) begin
      BtbPlugin_logic_memWrite_payload_mask = 1'b1;
    end
  end

  always @(*) begin
    BtbPlugin_logic_memWrite_payload_data_0_hash = BtbPlugin_logic_onLearn_hash;
    if(DecoderPlugin_logic_forgetPort_valid) begin
      BtbPlugin_logic_memWrite_payload_data_0_hash = (~ BtbPlugin_logic_onForget_hash);
    end
  end

  always @(*) begin
    BtbPlugin_logic_memWrite_payload_data_0_sliceLow = LearnPlugin_logic_learn_payload_pcOnLastSlice[1 : 1];
    if(DecoderPlugin_logic_forgetPort_valid) begin
      BtbPlugin_logic_memWrite_payload_data_0_sliceLow = DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice[1 : 1];
    end
  end

  assign BtbPlugin_logic_memWrite_payload_data_0_pcTarget = (LearnPlugin_logic_learn_payload_pcTarget >>> 1'd1);
  always @(*) begin
    BtbPlugin_logic_memWrite_payload_data_0_isBranch = LearnPlugin_logic_learn_payload_isBranch;
    if(DecoderPlugin_logic_forgetPort_valid) begin
      BtbPlugin_logic_memWrite_payload_data_0_isBranch = 1'b0;
    end
  end

  always @(*) begin
    BtbPlugin_logic_memWrite_payload_data_0_isPush = LearnPlugin_logic_learn_payload_isPush;
    if(DecoderPlugin_logic_forgetPort_valid) begin
      BtbPlugin_logic_memWrite_payload_data_0_isPush = 1'b0;
    end
  end

  always @(*) begin
    BtbPlugin_logic_memWrite_payload_data_0_isPop = LearnPlugin_logic_learn_payload_isPop;
    if(DecoderPlugin_logic_forgetPort_valid) begin
      BtbPlugin_logic_memWrite_payload_data_0_isPop = 1'b0;
    end
  end

  assign lane0_integer_WriteBackPlugin_logic_stages_0_hits = {lane0_IntFormatPlugin_logic_stages_0_wb_valid,early0_BranchPlugin_logic_wb_valid};
  assign lane0_integer_WriteBackPlugin_logic_stages_0_muxed = ((lane0_integer_WriteBackPlugin_logic_stages_0_hits[0] ? early0_BranchPlugin_logic_wb_payload : 64'h0) | (lane0_integer_WriteBackPlugin_logic_stages_0_hits[1] ? lane0_IntFormatPlugin_logic_stages_0_wb_payload : 64'h0));
  assign execute_ctrl2_lane0_integer_WriteBackPlugin_logic_DATA_lane0_bypass = lane0_integer_WriteBackPlugin_logic_stages_0_muxed;
  assign lane0_integer_WriteBackPlugin_logic_stages_0_write_valid = (((((execute_ctrl2_down_LANE_SEL_lane0 && execute_ctrl2_down_isReady) && (! execute_lane0_ctrls_2_downIsCancel)) && (|lane0_integer_WriteBackPlugin_logic_stages_0_hits)) && execute_ctrl2_up_RD_ENABLE_lane0) && execute_ctrl2_down_COMMIT_lane0);
  assign lane0_integer_WriteBackPlugin_logic_stages_0_write_payload_uopId = execute_ctrl2_down_Decode_UOP_ID_lane0;
  assign lane0_integer_WriteBackPlugin_logic_stages_0_write_payload_data = lane0_integer_WriteBackPlugin_logic_stages_0_muxed;
  assign lane0_integer_WriteBackPlugin_logic_stages_1_hits = lane0_IntFormatPlugin_logic_stages_2_wb_valid;
  assign lane0_integer_WriteBackPlugin_logic_stages_1_muxed = (lane0_integer_WriteBackPlugin_logic_stages_1_hits[0] ? lane0_IntFormatPlugin_logic_stages_2_wb_payload : 64'h0);
  assign lane0_integer_WriteBackPlugin_logic_stages_1_merged = (execute_ctrl3_up_lane0_integer_WriteBackPlugin_logic_DATA_lane0 | lane0_integer_WriteBackPlugin_logic_stages_1_muxed);
  assign execute_ctrl3_lane0_integer_WriteBackPlugin_logic_DATA_lane0_bypass = lane0_integer_WriteBackPlugin_logic_stages_1_merged;
  assign lane0_integer_WriteBackPlugin_logic_stages_1_write_valid = (((((execute_ctrl3_down_LANE_SEL_lane0 && execute_ctrl3_down_isReady) && (! execute_lane0_ctrls_3_downIsCancel)) && (|lane0_integer_WriteBackPlugin_logic_stages_1_hits)) && execute_ctrl3_up_RD_ENABLE_lane0) && execute_ctrl3_down_COMMIT_lane0);
  assign lane0_integer_WriteBackPlugin_logic_stages_1_write_payload_uopId = execute_ctrl3_down_Decode_UOP_ID_lane0;
  assign lane0_integer_WriteBackPlugin_logic_stages_1_write_payload_data = lane0_integer_WriteBackPlugin_logic_stages_1_muxed;
  assign lane0_integer_WriteBackPlugin_logic_stages_2_hits = lane0_IntFormatPlugin_logic_stages_1_wb_valid;
  assign lane0_integer_WriteBackPlugin_logic_stages_2_muxed = (lane0_integer_WriteBackPlugin_logic_stages_2_hits[0] ? lane0_IntFormatPlugin_logic_stages_1_wb_payload : 64'h0);
  assign lane0_integer_WriteBackPlugin_logic_stages_2_merged = (execute_ctrl4_up_lane0_integer_WriteBackPlugin_logic_DATA_lane0 | lane0_integer_WriteBackPlugin_logic_stages_2_muxed);
  assign execute_ctrl4_lane0_integer_WriteBackPlugin_logic_DATA_lane0_bypass = lane0_integer_WriteBackPlugin_logic_stages_2_merged;
  assign lane0_integer_WriteBackPlugin_logic_stages_2_write_valid = (((((execute_ctrl4_down_LANE_SEL_lane0 && execute_ctrl4_down_isReady) && (! execute_lane0_ctrls_4_downIsCancel)) && (|lane0_integer_WriteBackPlugin_logic_stages_2_hits)) && execute_ctrl4_up_RD_ENABLE_lane0) && execute_ctrl4_down_COMMIT_lane0);
  assign lane0_integer_WriteBackPlugin_logic_stages_2_write_payload_uopId = execute_ctrl4_down_Decode_UOP_ID_lane0;
  assign lane0_integer_WriteBackPlugin_logic_stages_2_write_payload_data = lane0_integer_WriteBackPlugin_logic_stages_2_muxed;
  assign lane0_integer_WriteBackPlugin_logic_write_port_valid = (((((execute_ctrl4_up_LANE_SEL_lane0 && execute_ctrl4_down_isReady) && (! execute_lane0_ctrls_4_upIsCancel)) && execute_ctrl4_up_RD_ENABLE_lane0) && execute_ctrl4_down_lane0_integer_WriteBackPlugin_SEL_lane0) && execute_ctrl4_down_COMMIT_lane0);
  assign lane0_integer_WriteBackPlugin_logic_write_port_address = execute_ctrl4_down_RD_PHYS_lane0[4 : 0];
  assign lane0_integer_WriteBackPlugin_logic_write_port_data = execute_ctrl4_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
  assign lane0_integer_WriteBackPlugin_logic_write_port_uopId = execute_ctrl4_down_Decode_UOP_ID_lane0;
  assign decode_ctrls_1_down_AguPlugin_CLEAN_0 = _zz_decode_ctrls_1_down_AguPlugin_CLEAN_0[0];
  assign decode_ctrls_1_down_AguPlugin_INVALIDATE_0 = _zz_decode_ctrls_1_down_AguPlugin_INVALIDATE_0[0];
  assign decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_0 = _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_0[0];
  assign decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_0 = _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_0[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0) == 32'h0);
  assign decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0[0];
  assign decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_0 = _zz_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_0[0];
  assign _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00002050) == 32'h00002050);
  assign _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_1 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00001050) == 32'h00001050);
  assign decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_0 = _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_0[0];
  assign decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_0 = _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_0[0];
  assign decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_0 = _zz_decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_0[0];
  assign decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_0 = _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_0[0];
  assign decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0 = _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_2[0];
  assign decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_0 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_0[0];
  assign decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0_1[0];
  assign when_CtrlLaneApi_l50_2 = (decode_ctrls_1_up_isReady || decode_ctrls_1_lane0_upIsCancel);
  assign WhiteboxerPlugin_logic_serializeds_0_fire = (decode_ctrls_1_up_LANE_SEL_0 && (! decode_ctrls_1_up_LANE_SEL_0_regNext_1));
  assign WhiteboxerPlugin_logic_serializeds_0_decodeId = decode_ctrls_1_down_Decode_DOP_ID_0;
  assign WhiteboxerPlugin_logic_serializeds_0_microOpId = decode_ctrls_1_down_Decode_UOP_ID_0;
  assign WhiteboxerPlugin_logic_serializeds_0_microOp = decode_ctrls_1_down_Decode_UOP_0;
  assign when_CtrlLaneApi_l50_3 = (execute_ctrl0_down_isReady || execute_lane0_ctrls_0_downIsCancel);
  assign WhiteboxerPlugin_logic_dispatches_0_fire = (execute_ctrl0_down_LANE_SEL_lane0 && (! execute_ctrl0_down_LANE_SEL_lane0_regNext));
  assign WhiteboxerPlugin_logic_dispatches_0_microOpId = execute_ctrl0_down_Decode_UOP_ID_lane0;
  assign when_CtrlLaneApi_l50_4 = (execute_ctrl2_down_isReady || execute_lane0_ctrls_2_downIsCancel);
  assign WhiteboxerPlugin_logic_executes_0_fire = ((execute_ctrl2_down_LANE_SEL_lane0 && (! execute_ctrl2_down_LANE_SEL_lane0_regNext)) && execute_ctrl2_down_COMMIT_lane0);
  assign WhiteboxerPlugin_logic_executes_0_microOpId = execute_ctrl2_down_Decode_UOP_ID_lane0;
  assign BtbPlugin_logic_onForget_hash = DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice[26 : 11];
  assign BtbPlugin_logic_memRead_cmd_valid = fetch_logic_ctrls_0_down_isReady;
  assign BtbPlugin_logic_memRead_cmd_payload = _zz_BtbPlugin_logic_memRead_cmd_payload[8:0];
  assign fetch_logic_ctrls_0_down_BtbPlugin_logic_readCmd_HAZARDS = ((BtbPlugin_logic_memWrite_valid && (BtbPlugin_logic_memWrite_payload_address == BtbPlugin_logic_memRead_cmd_payload)) ? BtbPlugin_logic_memWrite_payload_mask : 1'b0);
  assign fetch_logic_ctrls_0_haltRequest_BtbPlugin_l200 = BtbPlugin_logic_memWrite_valid;
  assign BtbPlugin_logic_predictions = {fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_1[1],fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0[1]};
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_hash = BtbPlugin_logic_memRead_rsp_0_hash;
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_sliceLow = BtbPlugin_logic_memRead_rsp_0_sliceLow;
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_pcTarget = BtbPlugin_logic_memRead_rsp_0_pcTarget;
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isBranch = BtbPlugin_logic_memRead_rsp_0_isBranch;
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isPush = BtbPlugin_logic_memRead_rsp_0_isPush;
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isPop = BtbPlugin_logic_memRead_rsp_0_isPop;
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_hitCalc_HIT = ((fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_hash == fetch_logic_ctrls_1_down_Fetch_WORD_PC[26 : 11]) && (fetch_logic_ctrls_1_down_Fetch_WORD_PC[1 : 1] <= fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_sliceLow));
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_predict_TAKEN = ((! fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isBranch) || BtbPlugin_logic_predictions[fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_sliceLow]);
  assign BtbPlugin_logic_ras_readIt = fetch_logic_ctrls_0_down_isReady;
  assign BtbPlugin_logic_applyIt_chunksMask = (fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_hitCalc_HIT && 1'b1);
  assign BtbPlugin_logic_applyIt_chunksTakenOh = (fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_predict_TAKEN & BtbPlugin_logic_applyIt_chunksMask);
  assign BtbPlugin_logic_applyIt_needIt = (fetch_logic_ctrls_1_up_isValid && (|BtbPlugin_logic_applyIt_chunksTakenOh));
  assign when_BtbPlugin_l233 = (fetch_logic_ctrls_1_up_isReady || fetch_logic_ctrls_1_up_isCancel);
  assign BtbPlugin_logic_applyIt_doIt = (BtbPlugin_logic_applyIt_needIt && (! BtbPlugin_logic_applyIt_correctionSent));
  assign BtbPlugin_logic_applyIt_entry_hash = fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_hash;
  assign BtbPlugin_logic_applyIt_entry_sliceLow = fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_sliceLow;
  assign BtbPlugin_logic_applyIt_entry_pcTarget = fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_pcTarget;
  assign BtbPlugin_logic_applyIt_entry_isBranch = fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isBranch;
  assign BtbPlugin_logic_applyIt_entry_isPush = fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isPush;
  assign BtbPlugin_logic_applyIt_entry_isPop = fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isPop;
  always @(*) begin
    BtbPlugin_logic_applyIt_pcTarget = BtbPlugin_logic_applyIt_entry_pcTarget;
    if(BtbPlugin_logic_applyIt_entry_isPop) begin
      BtbPlugin_logic_applyIt_pcTarget = BtbPlugin_logic_ras_read;
    end
  end

  assign BtbPlugin_logic_applyIt_doItSlice = BtbPlugin_logic_applyIt_entry_sliceLow;
  assign BtbPlugin_logic_applyIt_rasLogic_pushValid = (BtbPlugin_logic_applyIt_doIt && BtbPlugin_logic_applyIt_entry_isPush);
  always @(*) begin
    BtbPlugin_logic_applyIt_rasLogic_pushPc = fetch_logic_ctrls_1_down_Fetch_WORD_PC;
    BtbPlugin_logic_applyIt_rasLogic_pushPc[1 : 1] = BtbPlugin_logic_applyIt_doItSlice;
  end

  assign when_BtbPlugin_l246 = (BtbPlugin_logic_applyIt_doIt && BtbPlugin_logic_applyIt_entry_isPop);
  assign BtbPlugin_logic_flushPort_valid = BtbPlugin_logic_applyIt_doIt;
  assign BtbPlugin_logic_flushPort_payload_self = 1'b0;
  assign BtbPlugin_logic_pcPort_valid = BtbPlugin_logic_applyIt_doIt;
  assign BtbPlugin_logic_pcPort_payload_fault = 1'b0;
  assign BtbPlugin_logic_pcPort_payload_pc = ({1'd0,BtbPlugin_logic_applyIt_pcTarget} <<< 1'd1);
  assign fetch_logic_ctrls_1_down_Prediction_WORD_JUMPED = BtbPlugin_logic_applyIt_needIt;
  assign fetch_logic_ctrls_1_down_Prediction_WORD_JUMP_SLICE = BtbPlugin_logic_applyIt_doItSlice;
  assign fetch_logic_ctrls_1_down_Prediction_WORD_JUMP_PC = ({1'd0,BtbPlugin_logic_applyIt_pcTarget} <<< 1'd1);
  assign BtbPlugin_logic_applyIt_history_layers_0_history = fetch_logic_ctrls_1_down_Prediction_BRANCH_HISTORY;
  assign BtbPlugin_logic_applyIt_history_layersLogic_0_doIt = (BtbPlugin_logic_applyIt_chunksMask[0] && fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isBranch);
  assign BtbPlugin_logic_applyIt_history_layersLogic_0_shifted = {BtbPlugin_logic_applyIt_history_layers_0_history[10 : 0],fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_predict_TAKEN};
  assign BtbPlugin_logic_applyIt_history_layers_1_history = (BtbPlugin_logic_applyIt_history_layersLogic_0_doIt ? BtbPlugin_logic_applyIt_history_layersLogic_0_shifted : BtbPlugin_logic_applyIt_history_layers_0_history);
  assign BtbPlugin_logic_historyPort_valid = ((fetch_logic_ctrls_1_up_isValid && (! BtbPlugin_logic_applyIt_correctionSent)) && (|fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_hitCalc_HIT));
  assign BtbPlugin_logic_historyPort_payload_history = BtbPlugin_logic_applyIt_history_layers_1_history;
  always @(*) begin
    fetch_logic_ctrls_1_down_Prediction_WORD_SLICES_BRANCH[0] = ((fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_hitCalc_HIT && fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isBranch) && (fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_sliceLow == 1'b0));
    fetch_logic_ctrls_1_down_Prediction_WORD_SLICES_BRANCH[1] = ((fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_hitCalc_HIT && fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isBranch) && (fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_sliceLow == 1'b1));
  end

  always @(*) begin
    fetch_logic_ctrls_1_down_Prediction_WORD_SLICES_TAKEN[0] = fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_predict_TAKEN;
    fetch_logic_ctrls_1_down_Prediction_WORD_SLICES_TAKEN[1] = fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_predict_TAKEN;
  end

  assign AlignerPlugin_logic_buffer_flushIt = (|{(DecoderPlugin_logic_laneLogic_0_flushPort_valid && 1'b1),{(early0_EnvPlugin_logic_flushPort_valid && 1'b1),{(CsrAccessPlugin_logic_flushPort_valid && 1'b1),{(early0_BranchPlugin_logic_flushPort_valid && 1'b1),(LsuPlugin_logic_flushPort_valid && 1'b1)}}}});
  assign AlignerPlugin_logic_buffer_readers_0_firstFromBuffer = (|{_zz_AlignerPlugin_logic_extractors_0_redo_1,_zz_AlignerPlugin_logic_extractors_0_redo});
  assign AlignerPlugin_logic_buffer_readers_0_lastFromBuffer = ({AlignerPlugin_logic_extractors_0_usageMask[3],AlignerPlugin_logic_extractors_0_usageMask[2]} == 2'b00);
  assign _zz_AlignerPlugin_logic_extractors_0_ctx_instruction = {_zz_AlignerPlugin_logic_extractors_0_redo_3,{_zz_AlignerPlugin_logic_extractors_0_redo_2,{_zz_AlignerPlugin_logic_extractors_0_redo_1,_zz_AlignerPlugin_logic_extractors_0_redo}}};
  assign AlignerPlugin_logic_extractors_0_ctx_instruction = (((_zz_AlignerPlugin_logic_extractors_0_ctx_instruction[0] ? AlignerPlugin_logic_slicesInstructions_0 : 32'h0) | (_zz_AlignerPlugin_logic_extractors_0_ctx_instruction[1] ? AlignerPlugin_logic_slicesInstructions_1 : 32'h0)) | ((_zz_AlignerPlugin_logic_extractors_0_ctx_instruction[2] ? AlignerPlugin_logic_slicesInstructions_2 : 32'h0) | (_zz_AlignerPlugin_logic_extractors_0_ctx_instruction[3] ? AlignerPlugin_logic_slicesInstructions_3 : 32'h0)));
  always @(*) begin
    AlignerPlugin_logic_extractors_0_ctx_pc = (AlignerPlugin_logic_buffer_readers_0_firstFromBuffer ? AlignerPlugin_logic_buffer_pc : fetch_logic_ctrls_2_down_Fetch_WORD_PC);
    AlignerPlugin_logic_extractors_0_ctx_pc[1 : 1] = _zz_AlignerPlugin_logic_extractors_0_ctx_pc;
  end

  assign _zz_AlignerPlugin_logic_extractors_0_ctx_pc = (|{_zz_AlignerPlugin_logic_extractors_0_redo_3,_zz_AlignerPlugin_logic_extractors_0_redo_1});
  assign AlignerPlugin_logic_extractors_0_ctx_trap = ((AlignerPlugin_logic_buffer_readers_0_firstFromBuffer && AlignerPlugin_logic_buffer_trap) || ((! AlignerPlugin_logic_buffer_readers_0_lastFromBuffer) && fetch_logic_ctrls_2_down_TRAP));
  assign AlignerPlugin_logic_extractors_0_ctx_hm_Fetch_ID = (AlignerPlugin_logic_buffer_readers_0_firstFromBuffer ? AlignerPlugin_logic_buffer_hm_Fetch_ID : fetch_logic_ctrls_2_down_Fetch_ID);
  assign AlignerPlugin_logic_extractors_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_0 = (AlignerPlugin_logic_buffer_readers_0_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_GSharePlugin_GSHARE_COUNTER_0 : fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_0);
  assign AlignerPlugin_logic_extractors_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_1 = (AlignerPlugin_logic_buffer_readers_0_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_GSharePlugin_GSHARE_COUNTER_1 : fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_1);
  assign AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_BRANCH_HISTORY = (AlignerPlugin_logic_buffer_readers_0_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_Prediction_BRANCH_HISTORY : fetch_logic_ctrls_2_down_Prediction_BRANCH_HISTORY);
  assign AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_SLICES_BRANCH = (AlignerPlugin_logic_buffer_readers_0_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_Prediction_WORD_SLICES_BRANCH : fetch_logic_ctrls_2_down_Prediction_WORD_SLICES_BRANCH);
  assign AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_SLICES_TAKEN = (AlignerPlugin_logic_buffer_readers_0_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_Prediction_WORD_SLICES_TAKEN : fetch_logic_ctrls_2_down_Prediction_WORD_SLICES_TAKEN);
  assign AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_JUMP_PC = (AlignerPlugin_logic_buffer_readers_0_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_Prediction_WORD_JUMP_PC : fetch_logic_ctrls_2_down_Prediction_WORD_JUMP_PC);
  assign AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_JUMPED = (AlignerPlugin_logic_buffer_readers_0_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_Prediction_WORD_JUMPED : fetch_logic_ctrls_2_down_Prediction_WORD_JUMPED);
  assign AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_JUMP_SLICE = (AlignerPlugin_logic_buffer_readers_0_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_Prediction_WORD_JUMP_SLICE : fetch_logic_ctrls_2_down_Prediction_WORD_JUMP_SLICE);
  assign AlignerPlugin_api_downMoving = decode_ctrls_0_up_isMoving;
  always @(*) begin
    TrapPlugin_logic_harts_0_crsPorts_read_valid = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
        TrapPlugin_logic_harts_0_crsPorts_read_valid = 1'b1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_WAIT : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
        TrapPlugin_logic_harts_0_crsPorts_read_valid = 1'b1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_logic_harts_0_crsPorts_read_address = 4'bxxxx;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
        TrapPlugin_logic_harts_0_crsPorts_read_address = _zz_TrapPlugin_logic_harts_0_crsPorts_read_address;
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_WAIT : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
        TrapPlugin_logic_harts_0_crsPorts_read_address = _zz_TrapPlugin_logic_harts_0_crsPorts_read_address_1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  assign decode_logic_flushes_0_onLanes_0_doIt = (|{(DecoderPlugin_logic_laneLogic_0_flushPort_valid && 1'b1),{(early0_EnvPlugin_logic_flushPort_valid && 1'b1),{(CsrAccessPlugin_logic_flushPort_valid && 1'b1),{(early0_BranchPlugin_logic_flushPort_valid && 1'b1),(LsuPlugin_logic_flushPort_valid && 1'b1)}}}});
  assign decode_ctrls_0_lane0_downIsCancel = 1'b0;
  assign decode_ctrls_0_lane0_upIsCancel = decode_logic_flushes_0_onLanes_0_doIt;
  assign decode_logic_flushes_1_onLanes_0_doIt = (|{((DecoderPlugin_logic_laneLogic_0_flushPort_valid && 1'b1) && (1'b0 || (1'b1 && DecoderPlugin_logic_laneLogic_0_flushPort_payload_self))),{(early0_EnvPlugin_logic_flushPort_valid && 1'b1),{(CsrAccessPlugin_logic_flushPort_valid && 1'b1),{(early0_BranchPlugin_logic_flushPort_valid && 1'b1),(LsuPlugin_logic_flushPort_valid && 1'b1)}}}});
  assign decode_ctrls_1_lane0_downIsCancel = 1'b0;
  assign decode_ctrls_1_lane0_upIsCancel = decode_logic_flushes_1_onLanes_0_doIt;
  assign decode_logic_trapPending[0] = (|{((decode_ctrls_1_up_LANE_SEL_0 && 1'b1) && decode_ctrls_1_down_TRAP_0),((decode_ctrls_0_up_LANE_SEL_0 && 1'b1) && decode_ctrls_0_down_TRAP_0)});
  always @(*) begin
    TrapPlugin_logic_harts_0_crsPorts_write_valid = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
        TrapPlugin_logic_harts_0_crsPorts_write_valid = 1'b1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
        TrapPlugin_logic_harts_0_crsPorts_write_valid = 1'b1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_WAIT : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_logic_harts_0_crsPorts_write_address = 4'bxxxx;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
        TrapPlugin_logic_harts_0_crsPorts_write_address = _zz_TrapPlugin_logic_harts_0_crsPorts_write_address;
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
        TrapPlugin_logic_harts_0_crsPorts_write_address = _zz_TrapPlugin_logic_harts_0_crsPorts_write_address_1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_WAIT : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_logic_harts_0_crsPorts_write_data = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
        TrapPlugin_logic_harts_0_crsPorts_write_data = _zz_TrapPlugin_logic_harts_0_crsPorts_write_data;
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
        TrapPlugin_logic_harts_0_crsPorts_write_data = _zz_TrapPlugin_logic_harts_0_crsPorts_write_data_2;
        if(TrapPlugin_logic_harts_0_trap_fsm_triggerEbreakReg) begin
          TrapPlugin_logic_harts_0_crsPorts_write_data = _zz_TrapPlugin_logic_harts_0_crsPorts_write_data_4;
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_WAIT : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  assign TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_0_id = 4'b0001;
  assign TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_0_priority = 4'b0101;
  assign TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_0_privilege = 2'b01;
  assign TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_0_valid = ((_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_0_valid && (1'b1 && PrivilegedPlugin_logic_harts_0_m_ideleg_ss)) && (! 1'b0));
  assign TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_1_id = 4'b0101;
  assign TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_1_priority = 4'b0110;
  assign TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_1_privilege = 2'b01;
  assign TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_1_valid = ((_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_1_valid && (1'b1 && PrivilegedPlugin_logic_harts_0_m_ideleg_st)) && (! 1'b0));
  assign TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_2_id = 4'b1001;
  assign TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_2_priority = 4'b0100;
  assign TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_2_privilege = 2'b01;
  assign TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_2_valid = ((_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_2_valid && (1'b1 && PrivilegedPlugin_logic_harts_0_m_ideleg_se)) && (! 1'b0));
  assign _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_triggered_id = ((! TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_1_valid) || (TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_0_valid && ((TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_1_privilege < TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_0_privilege) || ((TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_0_privilege == TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_1_privilege) && (TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_0_priority < TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_1_priority)))));
  assign _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_triggered_priority = (_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_triggered_id ? TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_0_priority : TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_1_priority);
  assign _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_triggered_privilege = (_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_triggered_id ? TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_0_privilege : TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_1_privilege);
  assign _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_triggered_valid = (_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_triggered_id ? TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_0_valid : TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_1_valid);
  assign _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_triggered_id_1 = ((! TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_2_valid) || (_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_triggered_valid && ((TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_2_privilege < _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_triggered_privilege) || ((_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_triggered_privilege == TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_2_privilege) && (_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_triggered_priority < TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_2_priority)))));
  assign TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_0_id = 4'b0111;
  assign TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_0_priority = 4'b0011;
  assign TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_0_privilege = 2'b11;
  assign TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_0_valid = ((_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_0_valid && 1'b1) && (! 1'b0));
  assign TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_1_id = 4'b0011;
  assign TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_1_priority = 4'b0010;
  assign TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_1_privilege = 2'b11;
  assign TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_1_valid = ((_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_1_valid && 1'b1) && (! 1'b0));
  assign TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_2_id = 4'b1011;
  assign TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_2_priority = 4'b0001;
  assign TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_2_privilege = 2'b11;
  assign TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_2_valid = ((_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_2_valid && 1'b1) && (! 1'b0));
  assign TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_3_id = 4'b0001;
  assign TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_3_priority = 4'b0101;
  assign TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_3_privilege = 2'b11;
  assign TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_3_valid = ((_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_0_valid && 1'b1) && (! (|PrivilegedPlugin_logic_harts_0_m_ideleg_ss)));
  assign TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_4_id = 4'b0101;
  assign TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_4_priority = 4'b0110;
  assign TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_4_privilege = 2'b11;
  assign TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_4_valid = ((_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_1_valid && 1'b1) && (! (|PrivilegedPlugin_logic_harts_0_m_ideleg_st)));
  assign TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_5_id = 4'b1001;
  assign TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_5_priority = 4'b0100;
  assign TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_5_privilege = 2'b11;
  assign TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_5_valid = ((_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_2_valid && 1'b1) && (! (|PrivilegedPlugin_logic_harts_0_m_ideleg_se)));
  assign _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id = ((! TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_1_valid) || (TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_0_valid && ((TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_1_privilege < TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_0_privilege) || ((TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_0_privilege == TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_1_privilege) && (TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_0_priority < TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_1_priority)))));
  assign _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_1 = (_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id ? TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_0_priority : TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_1_priority);
  assign _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_2 = (_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id ? TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_0_privilege : TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_1_privilege);
  assign _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_3 = (_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id ? TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_0_valid : TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_1_valid);
  assign _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_4 = ((! TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_3_valid) || (TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_2_valid && ((TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_3_privilege < TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_2_privilege) || ((TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_2_privilege == TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_3_privilege) && (TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_2_priority < TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_3_priority)))));
  assign _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_5 = (_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_4 ? TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_2_priority : TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_3_priority);
  assign _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_6 = (_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_4 ? TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_2_privilege : TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_3_privilege);
  assign _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_7 = (_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_4 ? TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_2_valid : TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_3_valid);
  assign _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_8 = ((! TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_5_valid) || (TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_4_valid && ((TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_5_privilege < TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_4_privilege) || ((TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_4_privilege == TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_5_privilege) && (TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_4_priority < TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_5_priority)))));
  assign _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_priority = (_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_8 ? TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_4_priority : TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_5_priority);
  assign _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_privilege = (_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_8 ? TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_4_privilege : TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_5_privilege);
  assign _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_valid = (_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_8 ? TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_4_valid : TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_5_valid);
  assign _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_9 = ((! _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_7) || (_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_3 && ((_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_6 < _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_2) || ((_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_2 == _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_6) && (_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_1 < _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_5)))));
  assign _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_priority_1 = (_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_9 ? _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_1 : _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_5);
  assign _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_privilege_1 = (_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_9 ? _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_2 : _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_6);
  assign _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_valid_1 = (_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_9 ? _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_3 : _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_7);
  assign _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_10 = ((! _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_valid) || (_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_valid_1 && ((_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_privilege < _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_privilege_1) || ((_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_privilege_1 == _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_privilege) && (_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_priority_1 < _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_priority)))));
  assign TrapPlugin_logic_harts_0_interrupt_xtopi_0_int = (TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_triggered_valid ? TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_triggered_id : 4'b0000);
  assign TrapPlugin_logic_harts_0_interrupt_xtopi_1_int = (TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_valid ? TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id : 4'b0000);
  assign _zz_TrapPlugin_logic_harts_0_interrupt_result_privilege = TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_triggered_privilege;
  assign _zz_TrapPlugin_logic_harts_0_interrupt_result_valid = (TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_triggered_valid && ((PrivilegedPlugin_logic_harts_0_s_status_sie && (! PrivilegedPlugin_logic_harts_0_withMachinePrivilege)) || (! PrivilegedPlugin_logic_harts_0_withSupervisorPrivilege)));
  assign _zz_TrapPlugin_logic_harts_0_interrupt_result_privilege_1 = TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_privilege;
  assign _zz_TrapPlugin_logic_harts_0_interrupt_result_valid_1 = (TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_valid && (PrivilegedPlugin_logic_harts_0_m_status_mie || (! PrivilegedPlugin_logic_harts_0_withMachinePrivilege)));
  assign _zz_TrapPlugin_logic_harts_0_interrupt_result_id = ((! _zz_TrapPlugin_logic_harts_0_interrupt_result_valid_1) || (_zz_TrapPlugin_logic_harts_0_interrupt_result_valid && (_zz_TrapPlugin_logic_harts_0_interrupt_result_privilege_1 < _zz_TrapPlugin_logic_harts_0_interrupt_result_privilege)));
  assign TrapPlugin_logic_harts_0_interrupt_result_id = (_zz_TrapPlugin_logic_harts_0_interrupt_result_id ? TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_triggered_id : TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id);
  assign TrapPlugin_logic_harts_0_interrupt_result_priority = (_zz_TrapPlugin_logic_harts_0_interrupt_result_id ? TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_triggered_priority : TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_priority);
  assign TrapPlugin_logic_harts_0_interrupt_result_privilege = (_zz_TrapPlugin_logic_harts_0_interrupt_result_id ? _zz_TrapPlugin_logic_harts_0_interrupt_result_privilege : _zz_TrapPlugin_logic_harts_0_interrupt_result_privilege_1);
  assign TrapPlugin_logic_harts_0_interrupt_result_valid = (_zz_TrapPlugin_logic_harts_0_interrupt_result_id ? _zz_TrapPlugin_logic_harts_0_interrupt_result_valid : _zz_TrapPlugin_logic_harts_0_interrupt_result_valid_1);
  assign TrapPlugin_logic_harts_0_interrupt_valid = TrapPlugin_logic_harts_0_interrupt_result_valid;
  assign TrapPlugin_logic_harts_0_interrupt_code = TrapPlugin_logic_harts_0_interrupt_result_id;
  assign TrapPlugin_logic_harts_0_interrupt_targetPrivilege = TrapPlugin_logic_harts_0_interrupt_result_privilege;
  assign TrapPlugin_logic_harts_0_interrupt_pendingInterrupt = (TrapPlugin_logic_harts_0_interrupt_validBuffer && PrivilegedPlugin_api_harts_0_allowInterrupts);
  assign when_TrapPlugin_l269 = (|{_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_2_valid,{_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_1_valid,{_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_0_valid,{_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_2_valid,{_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_1_valid,_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_0_valid}}}}});
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid = (early0_EnvPlugin_logic_trapPort_valid && 1'b1);
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_valid = (FetchL1Plugin_logic_trapPort_valid && 1'b1);
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_valid = (LsuPlugin_logic_trapPort_valid && 1'b1);
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid_1 = (CsrAccessPlugin_logic_trapPort_valid && 1'b1);
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid = (DecoderPlugin_logic_laneLogic_0_trapPort_valid && 1'b1);
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_valid = (|_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_valid);
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_exception = LsuPlugin_logic_trapPort_payload_exception;
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_tval = LsuPlugin_logic_trapPort_payload_tval;
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_code = LsuPlugin_logic_trapPort_payload_code;
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_arg = LsuPlugin_logic_trapPort_payload_arg;
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_exception = {(_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid_1 && (&(! (_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid && 1'b0)))),(_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid && (&(! (_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid_1 && 1'b0))))};
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid = (|{_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid_1,_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid});
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_exception_1 = ((_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_exception[0] ? {early0_EnvPlugin_logic_trapPort_payload_arg,{early0_EnvPlugin_logic_trapPort_payload_code,{early0_EnvPlugin_logic_trapPort_payload_tval,early0_EnvPlugin_logic_trapPort_payload_exception}}} : 47'h0) | (_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_exception[1] ? {CsrAccessPlugin_logic_trapPort_payload_arg,{CsrAccessPlugin_logic_trapPort_payload_code,{CsrAccessPlugin_logic_trapPort_payload_tval,CsrAccessPlugin_logic_trapPort_payload_exception}}} : 47'h0));
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_exception = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_exception_1[0];
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_tval = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_exception_1[39 : 1];
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_code = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_exception_1[43 : 40];
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_arg = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_exception_1[46 : 44];
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid = (|_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid);
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_exception = DecoderPlugin_logic_laneLogic_0_trapPort_payload_exception;
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_tval = DecoderPlugin_logic_laneLogic_0_trapPort_payload_tval;
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_code = DecoderPlugin_logic_laneLogic_0_trapPort_payload_code;
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_arg = DecoderPlugin_logic_laneLogic_0_trapPort_payload_arg;
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_valid = (|_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_valid);
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_exception = FetchL1Plugin_logic_trapPort_payload_exception;
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_tval = FetchL1Plugin_logic_trapPort_payload_tval;
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_code = FetchL1Plugin_logic_trapPort_payload_code;
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_arg = FetchL1Plugin_logic_trapPort_payload_arg;
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh = {TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_valid,{TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid,{TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid,TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_valid}}};
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_1 = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh[0];
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_2 = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh[1];
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_3 = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh[2];
  always @(*) begin
    _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_4[0] = (_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_1 && (! 1'b0));
    _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_4[1] = (_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_2 && (! _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_1));
    _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_4[2] = (_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_3 && (! (|{_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_2,_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_1})));
    _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_4[3] = (_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh[3] && (! (|{_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_3,{_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_2,_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_1}})));
  end

  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_oh = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_4;
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_down_valid = (|{_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid,{_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid_1,{_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_valid,{_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_valid,_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid}}}});
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception = (((TrapPlugin_logic_harts_0_trap_pending_arbiter_oh[0] ? {TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_arg,{TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_code,_zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception}} : 47'h0) | (TrapPlugin_logic_harts_0_trap_pending_arbiter_oh[1] ? {TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_arg,{TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_code,_zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception_1}} : 47'h0)) | ((TrapPlugin_logic_harts_0_trap_pending_arbiter_oh[2] ? {TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_arg,{TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_code,_zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception_2}} : 47'h0) | (TrapPlugin_logic_harts_0_trap_pending_arbiter_oh[3] ? {TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_arg,{TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_code,_zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception_3}} : 47'h0)));
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception[0];
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_tval = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception[39 : 1];
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_code = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception[43 : 40];
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_arg = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception[46 : 44];
  assign TrapPlugin_logic_harts_0_trap_pending_xret_sourcePrivilege = TrapPlugin_logic_harts_0_trap_pending_state_arg[1 : 0];
  always @(*) begin
    TrapPlugin_logic_harts_0_trap_pending_xret_targetPrivilege = PrivilegedPlugin_logic_harts_0_m_status_mpp;
    case(TrapPlugin_logic_harts_0_trap_pending_xret_sourcePrivilege)
      2'b01 : begin
        TrapPlugin_logic_harts_0_trap_pending_xret_targetPrivilege = {1'b0,PrivilegedPlugin_logic_harts_0_s_status_spp};
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_logic_harts_0_trap_exception_exceptionTargetPrivilegeUncapped = 2'b11;
    case(TrapPlugin_logic_harts_0_trap_exception_code)
      4'b0000 : begin
        if(when_TrapPlugin_l306) begin
          TrapPlugin_logic_harts_0_trap_exception_exceptionTargetPrivilegeUncapped = 2'b01;
        end
      end
      4'b0011 : begin
        if(when_TrapPlugin_l306_1) begin
          TrapPlugin_logic_harts_0_trap_exception_exceptionTargetPrivilegeUncapped = 2'b01;
        end
      end
      4'b1000 : begin
        if(when_TrapPlugin_l306_2) begin
          TrapPlugin_logic_harts_0_trap_exception_exceptionTargetPrivilegeUncapped = 2'b01;
        end
      end
      4'b1001 : begin
        if(when_TrapPlugin_l306_3) begin
          TrapPlugin_logic_harts_0_trap_exception_exceptionTargetPrivilegeUncapped = 2'b01;
        end
      end
      4'b1100 : begin
        if(when_TrapPlugin_l306_4) begin
          TrapPlugin_logic_harts_0_trap_exception_exceptionTargetPrivilegeUncapped = 2'b01;
        end
      end
      4'b1101 : begin
        if(when_TrapPlugin_l306_5) begin
          TrapPlugin_logic_harts_0_trap_exception_exceptionTargetPrivilegeUncapped = 2'b01;
        end
      end
      4'b1111 : begin
        if(when_TrapPlugin_l306_6) begin
          TrapPlugin_logic_harts_0_trap_exception_exceptionTargetPrivilegeUncapped = 2'b01;
        end
      end
      default : begin
      end
    endcase
  end

  assign TrapPlugin_logic_harts_0_trap_exception_code = TrapPlugin_logic_harts_0_trap_pending_state_code;
  assign when_TrapPlugin_l306 = ((1'b1 && PrivilegedPlugin_logic_harts_0_m_edeleg_iam) && (! 1'b0));
  assign when_TrapPlugin_l306_1 = ((1'b1 && PrivilegedPlugin_logic_harts_0_m_edeleg_bp) && (! 1'b0));
  assign when_TrapPlugin_l306_2 = ((1'b1 && PrivilegedPlugin_logic_harts_0_m_edeleg_eu) && (! 1'b0));
  assign when_TrapPlugin_l306_3 = ((1'b1 && PrivilegedPlugin_logic_harts_0_m_edeleg_es) && (! 1'b0));
  assign when_TrapPlugin_l306_4 = ((1'b1 && PrivilegedPlugin_logic_harts_0_m_edeleg_ipf) && (! 1'b0));
  assign when_TrapPlugin_l306_5 = ((1'b1 && PrivilegedPlugin_logic_harts_0_m_edeleg_lpf) && (! 1'b0));
  assign when_TrapPlugin_l306_6 = ((1'b1 && PrivilegedPlugin_logic_harts_0_m_edeleg_spf) && (! 1'b0));
  assign TrapPlugin_logic_harts_0_trap_exception_targetPrivilege = ((PrivilegedPlugin_logic_harts_0_privilege < TrapPlugin_logic_harts_0_trap_exception_exceptionTargetPrivilegeUncapped) ? TrapPlugin_logic_harts_0_trap_exception_exceptionTargetPrivilegeUncapped : PrivilegedPlugin_logic_harts_0_privilege);
  assign PrivilegedPlugin_logic_harts_0_commitMask = (((execute_ctrl5_down_LANE_SEL_lane0 && execute_ctrl5_down_isReady) && (! execute_lane0_ctrls_5_downIsCancel)) && execute_ctrl5_down_COMMIT_lane0);
  assign TrapPlugin_logic_harts_0_trap_trigger_oh = (((execute_ctrl4_down_LANE_SEL_lane0 && execute_ctrl4_down_isReady) && (! execute_lane0_ctrls_4_downIsCancel)) && execute_ctrl4_down_TRAP_lane0);
  assign TrapPlugin_logic_harts_0_trap_trigger_valid = (|TrapPlugin_logic_harts_0_trap_trigger_oh);
  always @(*) begin
    TrapPlugin_logic_harts_0_trap_whitebox_trap = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_WAIT : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
        TrapPlugin_logic_harts_0_trap_whitebox_trap = 1'b1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_logic_harts_0_trap_whitebox_interrupt = 1'bx;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_WAIT : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
        TrapPlugin_logic_harts_0_trap_whitebox_interrupt = TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_interrupt;
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_logic_harts_0_trap_whitebox_code = 4'bxxxx;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_WAIT : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
        TrapPlugin_logic_harts_0_trap_whitebox_code = TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_code;
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_logic_harts_0_trap_historyPort_valid = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
        TrapPlugin_logic_harts_0_trap_historyPort_valid = 1'b1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_WAIT : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  assign TrapPlugin_logic_harts_0_trap_historyPort_payload_history = TrapPlugin_logic_harts_0_trap_pending_history;
  always @(*) begin
    TrapPlugin_logic_harts_0_trap_pcPort_valid = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
        if(!when_TrapPlugin_l453) begin
          case(TrapPlugin_logic_harts_0_trap_pending_state_code)
            4'b0000 : begin
              TrapPlugin_logic_harts_0_trap_pcPort_valid = 1'b1;
            end
            4'b0001 : begin
            end
            4'b0010 : begin
            end
            4'b0100 : begin
            end
            4'b0101 : begin
            end
            4'b1000 : begin
            end
            4'b0110 : begin
            end
            4'b0111 : begin
            end
            default : begin
            end
          endcase
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_WAIT : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
        TrapPlugin_logic_harts_0_trap_pcPort_valid = 1'b1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
        TrapPlugin_logic_harts_0_trap_pcPort_valid = 1'b1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
        TrapPlugin_logic_harts_0_trap_pcPort_valid = 1'b1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  assign TrapPlugin_logic_harts_0_trap_pcPort_payload_fault = 1'b0;
  always @(*) begin
    TrapPlugin_logic_harts_0_trap_pcPort_payload_pc = 39'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
        if(!when_TrapPlugin_l453) begin
          case(TrapPlugin_logic_harts_0_trap_pending_state_code)
            4'b0000 : begin
              TrapPlugin_logic_harts_0_trap_pcPort_payload_pc = TrapPlugin_logic_harts_0_trap_pending_pc;
            end
            4'b0001 : begin
            end
            4'b0010 : begin
            end
            4'b0100 : begin
            end
            4'b0101 : begin
            end
            4'b1000 : begin
            end
            4'b0110 : begin
            end
            4'b0111 : begin
            end
            default : begin
            end
          endcase
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_WAIT : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
        TrapPlugin_logic_harts_0_trap_pcPort_payload_pc = _zz_TrapPlugin_logic_harts_0_trap_pcPort_payload_pc[38:0];
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
        TrapPlugin_logic_harts_0_trap_pcPort_payload_pc = _zz_TrapPlugin_logic_harts_0_trap_pcPort_payload_pc_1[38:0];
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
        TrapPlugin_logic_harts_0_trap_pcPort_payload_pc = TrapPlugin_logic_harts_0_trap_fsm_jumpTarget;
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  assign TrapPlugin_logic_harts_0_trap_fsm_wantExit = 1'b0;
  always @(*) begin
    TrapPlugin_logic_harts_0_trap_fsm_wantStart = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_WAIT : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
        TrapPlugin_logic_harts_0_trap_fsm_wantStart = 1'b1;
      end
    endcase
  end

  assign TrapPlugin_logic_harts_0_trap_fsm_wantKill = 1'b0;
  assign TrapPlugin_logic_harts_0_trap_fsm_inflightTrap = (|{execute_lane0_logic_trapPending[0],{DispatchPlugin_logic_trapPendings[0],decode_logic_trapPending[0]}});
  assign TrapPlugin_logic_harts_0_trap_fsm_holdPort = (TrapPlugin_logic_harts_0_trap_fsm_inflightTrap || (! (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_RUNNING)));
  assign TrapPlugin_api_harts_0_fsmBusy = (! (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_RUNNING));
  always @(*) begin
    TrapPlugin_logic_harts_0_trap_fsm_wfi = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
        if(!when_TrapPlugin_l453) begin
          case(TrapPlugin_logic_harts_0_trap_pending_state_code)
            4'b0000 : begin
            end
            4'b0001 : begin
            end
            4'b0010 : begin
            end
            4'b0100 : begin
            end
            4'b0101 : begin
            end
            4'b1000 : begin
              TrapPlugin_logic_harts_0_trap_fsm_wfi = 1'b1;
            end
            4'b0110 : begin
            end
            4'b0111 : begin
            end
            default : begin
            end
          endcase
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_WAIT : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_logic_harts_0_trap_fsm_buffer_sampleIt = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
        if(TrapPlugin_logic_harts_0_trap_trigger_valid) begin
          TrapPlugin_logic_harts_0_trap_fsm_buffer_sampleIt = 1'b1;
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_WAIT : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  assign TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_interrupt = ((TrapPlugin_logic_harts_0_trap_pending_state_code == 4'b0000) && TrapPlugin_logic_harts_0_trap_fsm_buffer_i_valid);
  assign TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_targetPrivilege = (TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_interrupt ? TrapPlugin_logic_harts_0_trap_fsm_buffer_i_targetPrivilege : TrapPlugin_logic_harts_0_trap_exception_targetPrivilege);
  assign TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_tval = ((! TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_interrupt) ? TrapPlugin_logic_harts_0_trap_pending_state_tval : 39'h0);
  assign TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_code = (TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_interrupt ? TrapPlugin_logic_harts_0_trap_fsm_buffer_i_code : TrapPlugin_logic_harts_0_trap_pending_state_code);
  assign TrapPlugin_logic_harts_0_trap_fsm_resetToRunConditions_0 = (! TrapPlugin_logic_initHold);
  always @(*) begin
    TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_cmd_valid = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
        if(!when_TrapPlugin_l453) begin
          case(TrapPlugin_logic_harts_0_trap_pending_state_code)
            4'b0000 : begin
            end
            4'b0001 : begin
            end
            4'b0010 : begin
            end
            4'b0100 : begin
            end
            4'b0101 : begin
            end
            4'b1000 : begin
            end
            4'b0110 : begin
            end
            4'b0111 : begin
              TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_cmd_valid = 1'b1;
            end
            default : begin
            end
          endcase
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_WAIT : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  assign bits_storageEnable = 1'b1;
  assign bits_address = TrapPlugin_logic_harts_0_trap_pending_state_tval;
  assign bits_storageId = TrapPlugin_logic_harts_0_trap_pending_state_arg[2 : 2];
  always @(*) begin
    TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidate_cmd_valid = 1'b0;
    if(when_TrapPlugin_l399) begin
      TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidate_cmd_valid = 1'b1;
    end
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
        if(!when_TrapPlugin_l453) begin
          case(TrapPlugin_logic_harts_0_trap_pending_state_code)
            4'b0000 : begin
            end
            4'b0001 : begin
            end
            4'b0010 : begin
            end
            4'b0100 : begin
            end
            4'b0101 : begin
            end
            4'b1000 : begin
            end
            4'b0110 : begin
              TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidate_cmd_valid = 1'b1;
            end
            4'b0111 : begin
            end
            default : begin
            end
          endcase
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_WAIT : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  assign TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidate_cmd_fire = (TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidate_cmd_valid && TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidate_cmd_ready);
  assign when_TrapPlugin_l399 = (! TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidated);
  assign TrapPlugin_logic_harts_0_trap_fsm_jumpOffset = ((|{(TrapPlugin_logic_harts_0_trap_pending_state_code == 4'b1000),{(TrapPlugin_logic_harts_0_trap_pending_state_code == 4'b0110),{(TrapPlugin_logic_harts_0_trap_pending_state_code == 4'b0010),(TrapPlugin_logic_harts_0_trap_pending_state_code == 4'b0101)}}}) ? TrapPlugin_logic_harts_0_trap_pending_slices : 2'b00);
  always @(*) begin
    TrapPlugin_logic_fetchL1Invalidate_0_cmd_valid = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_WAIT : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
        TrapPlugin_logic_fetchL1Invalidate_0_cmd_valid = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_logic_lsuL1Invalidate_0_cmd_valid = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_WAIT : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
        TrapPlugin_logic_lsuL1Invalidate_0_cmd_valid = 1'b1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  assign TrapPlugin_logic_harts_0_trap_fsm_triggerEbreak = 1'b0;
  assign when_TrapPlugin_l602 = (TrapPlugin_logic_harts_0_crsPorts_read_valid && TrapPlugin_logic_harts_0_crsPorts_read_ready);
  assign TrapPlugin_logic_harts_0_trap_fsm_xretPrivilege = TrapPlugin_logic_harts_0_trap_pending_state_arg[1 : 0];
  assign PcPlugin_logic_forcedSpawn = (|{TrapPlugin_logic_harts_0_trap_pcPort_valid,{early0_BranchPlugin_logic_pcPort_valid,BtbPlugin_logic_pcPort_valid}});
  assign PcPlugin_logic_harts_0_self_pc = (PcPlugin_logic_harts_0_self_state + _zz_PcPlugin_logic_harts_0_self_pc);
  assign PcPlugin_logic_harts_0_self_flow_valid = 1'b1;
  assign PcPlugin_logic_harts_0_self_flow_payload_fault = PcPlugin_logic_harts_0_self_fault;
  assign PcPlugin_logic_harts_0_self_flow_payload_pc = PcPlugin_logic_harts_0_self_pc;
  assign PcPlugin_logic_harts_0_aggregator_sortedByPriority_2_laneValid = 1'b1;
  assign PcPlugin_logic_harts_0_aggregator_sortedByPriority_1_laneValid = 1'b1;
  assign PcPlugin_logic_harts_0_aggregator_sortedByPriority_0_laneValid = 1'b1;
  assign PcPlugin_logic_harts_0_aggregator_sortedByPriority_3_laneValid = 1'b1;
  assign PcPlugin_logic_harts_0_aggregator_valids_0 = ((TrapPlugin_logic_harts_0_trap_pcPort_valid && 1'b1) && PcPlugin_logic_harts_0_aggregator_sortedByPriority_0_laneValid);
  assign PcPlugin_logic_harts_0_aggregator_valids_1 = ((early0_BranchPlugin_logic_pcPort_valid && 1'b1) && PcPlugin_logic_harts_0_aggregator_sortedByPriority_1_laneValid);
  assign PcPlugin_logic_harts_0_aggregator_valids_2 = ((BtbPlugin_logic_pcPort_valid && 1'b1) && PcPlugin_logic_harts_0_aggregator_sortedByPriority_2_laneValid);
  assign PcPlugin_logic_harts_0_aggregator_valids_3 = ((PcPlugin_logic_harts_0_self_flow_valid && 1'b1) && PcPlugin_logic_harts_0_aggregator_sortedByPriority_3_laneValid);
  assign _zz_PcPlugin_logic_harts_0_aggregator_oh = {PcPlugin_logic_harts_0_aggregator_valids_3,{PcPlugin_logic_harts_0_aggregator_valids_2,{PcPlugin_logic_harts_0_aggregator_valids_1,PcPlugin_logic_harts_0_aggregator_valids_0}}};
  assign _zz_PcPlugin_logic_harts_0_aggregator_oh_1 = _zz_PcPlugin_logic_harts_0_aggregator_oh[0];
  assign _zz_PcPlugin_logic_harts_0_aggregator_oh_2 = _zz_PcPlugin_logic_harts_0_aggregator_oh[1];
  assign _zz_PcPlugin_logic_harts_0_aggregator_oh_3 = _zz_PcPlugin_logic_harts_0_aggregator_oh[2];
  always @(*) begin
    _zz_PcPlugin_logic_harts_0_aggregator_oh_4[0] = (_zz_PcPlugin_logic_harts_0_aggregator_oh_1 && (! 1'b0));
    _zz_PcPlugin_logic_harts_0_aggregator_oh_4[1] = (_zz_PcPlugin_logic_harts_0_aggregator_oh_2 && (! _zz_PcPlugin_logic_harts_0_aggregator_oh_1));
    _zz_PcPlugin_logic_harts_0_aggregator_oh_4[2] = (_zz_PcPlugin_logic_harts_0_aggregator_oh_3 && (! (|{_zz_PcPlugin_logic_harts_0_aggregator_oh_2,_zz_PcPlugin_logic_harts_0_aggregator_oh_1})));
    _zz_PcPlugin_logic_harts_0_aggregator_oh_4[3] = (_zz_PcPlugin_logic_harts_0_aggregator_oh[3] && (! (|{_zz_PcPlugin_logic_harts_0_aggregator_oh_3,{_zz_PcPlugin_logic_harts_0_aggregator_oh_2,_zz_PcPlugin_logic_harts_0_aggregator_oh_1}})));
  end

  assign PcPlugin_logic_harts_0_aggregator_oh = _zz_PcPlugin_logic_harts_0_aggregator_oh_4;
  assign _zz_PcPlugin_logic_harts_0_aggregator_target = PcPlugin_logic_harts_0_aggregator_oh[0];
  assign _zz_PcPlugin_logic_harts_0_aggregator_target_1 = PcPlugin_logic_harts_0_aggregator_oh[1];
  assign _zz_PcPlugin_logic_harts_0_aggregator_target_2 = PcPlugin_logic_harts_0_aggregator_oh[3];
  assign PcPlugin_logic_harts_0_aggregator_target = (((_zz_PcPlugin_logic_harts_0_aggregator_target ? TrapPlugin_logic_harts_0_trap_pcPort_payload_pc : 39'h0) | (_zz_PcPlugin_logic_harts_0_aggregator_target_1 ? early0_BranchPlugin_logic_pcPort_payload_pc : 39'h0)) | (_zz_PcPlugin_logic_harts_0_aggregator_target_2 ? PcPlugin_logic_harts_0_self_flow_payload_pc : 39'h0));
  assign PcPlugin_logic_harts_0_aggregator_fault = _zz_PcPlugin_logic_harts_0_aggregator_fault[0];
  assign _zz_PcPlugin_logic_harts_0_aggregator_fault_1 = PcPlugin_logic_harts_0_aggregator_oh[2];
  assign when_PcPlugin_l80 = (|_zz_PcPlugin_logic_harts_0_aggregator_fault_1);
  assign PcPlugin_logic_harts_0_holdComb = (|TrapPlugin_logic_harts_0_trap_fsm_holdPort);
  assign PcPlugin_logic_harts_0_output_valid = (! PcPlugin_logic_harts_0_holdReg);
  assign PcPlugin_logic_harts_0_output_payload_fault = PcPlugin_logic_harts_0_aggregator_fault_1;
  always @(*) begin
    PcPlugin_logic_harts_0_output_payload_pc = PcPlugin_logic_harts_0_aggregator_target_1;
    PcPlugin_logic_harts_0_output_payload_pc[0 : 0] = 1'b0;
  end

  assign PcPlugin_logic_harts_0_output_fire = (PcPlugin_logic_harts_0_output_valid && PcPlugin_logic_harts_0_output_ready);
  assign fetch_logic_ctrls_0_up_valid = PcPlugin_logic_harts_0_output_valid;
  assign PcPlugin_logic_harts_0_output_ready = fetch_logic_ctrls_0_up_ready;
  assign fetch_logic_ctrls_0_up_Fetch_WORD_PC = PcPlugin_logic_harts_0_output_payload_pc;
  assign fetch_logic_ctrls_0_up_Fetch_PC_FAULT = PcPlugin_logic_harts_0_output_payload_fault;
  always @(*) begin
    fetch_logic_ctrls_0_up_Fetch_ID = 10'bxxxxxxxxxx;
    fetch_logic_ctrls_0_up_Fetch_ID = PcPlugin_logic_harts_0_self_id;
  end

  assign PcPlugin_logic_holdHalter_doIt = PcPlugin_logic_harts_0_holdComb;
  assign fetch_logic_ctrls_0_haltRequest_PcPlugin_l133 = PcPlugin_logic_holdHalter_doIt;
  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_0_write_mask = 2'b00;
    if(!when_MmuPlugin_l565) begin
      FetchL1Plugin_logic_translationStorage_logic_sl_0_write_mask = 2'b11;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
        FetchL1Plugin_logic_translationStorage_logic_sl_0_write_mask = (MmuPlugin_logic_refill_storageOhReg[0] ? _zz_FetchL1Plugin_logic_translationStorage_logic_sl_0_write_mask : 2'b00);
        if(when_MmuPlugin_l505) begin
          FetchL1Plugin_logic_translationStorage_logic_sl_0_write_mask = 2'b00;
        end
      end
      MmuPlugin_logic_refill_DONE_1 : begin
      end
      MmuPlugin_logic_refill_DONE_2 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_0_write_address = 5'bxxxxx;
    if(!when_MmuPlugin_l565) begin
      FetchL1Plugin_logic_translationStorage_logic_sl_0_write_address = MmuPlugin_logic_invalidate_counter;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
        FetchL1Plugin_logic_translationStorage_logic_sl_0_write_address = MmuPlugin_logic_refill_virtual[16 : 12];
      end
      MmuPlugin_logic_refill_DONE_1 : begin
      end
      MmuPlugin_logic_refill_DONE_2 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_valid = 1'bx;
    if(!when_MmuPlugin_l565) begin
      FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_valid = 1'b0;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
        FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_valid = 1'b1;
      end
      MmuPlugin_logic_refill_DONE_1 : begin
      end
      MmuPlugin_logic_refill_DONE_2 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_virtualAddress = 22'bxxxxxxxxxxxxxxxxxxxxxx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
        FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_virtualAddress = MmuPlugin_logic_refill_virtual[38 : 17];
      end
      MmuPlugin_logic_refill_DONE_1 : begin
      end
      MmuPlugin_logic_refill_DONE_2 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_physicalAddress = 20'bxxxxxxxxxxxxxxxxxxxx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
        FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_physicalAddress = _zz_FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_physicalAddress[19:0];
      end
      MmuPlugin_logic_refill_DONE_1 : begin
      end
      MmuPlugin_logic_refill_DONE_2 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowRead = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
        FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowRead = MmuPlugin_logic_refill_load_flags_R;
      end
      MmuPlugin_logic_refill_DONE_1 : begin
      end
      MmuPlugin_logic_refill_DONE_2 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowWrite = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
        FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowWrite = (MmuPlugin_logic_refill_load_flags_W && MmuPlugin_logic_refill_load_flags_D);
      end
      MmuPlugin_logic_refill_DONE_1 : begin
      end
      MmuPlugin_logic_refill_DONE_2 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowExecute = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
        FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowExecute = MmuPlugin_logic_refill_load_flags_X;
      end
      MmuPlugin_logic_refill_DONE_1 : begin
      end
      MmuPlugin_logic_refill_DONE_2 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowUser = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
        FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowUser = MmuPlugin_logic_refill_load_flags_U;
      end
      MmuPlugin_logic_refill_DONE_1 : begin
      end
      MmuPlugin_logic_refill_DONE_2 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_willIncrement = 1'b0;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
        if(!when_MmuPlugin_l505) begin
          FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_willIncrement = 1'b1;
        end
      end
      MmuPlugin_logic_refill_DONE_1 : begin
      end
      MmuPlugin_logic_refill_DONE_2 : begin
      end
      default : begin
      end
    endcase
  end

  assign FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_willClear = 1'b0;
  assign FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_willOverflowIfInc = (FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_value == 1'b1);
  assign FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_willOverflow = (FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_willOverflowIfInc && FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_willIncrement);
  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_valueNext = (FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_value + FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_willIncrement);
    if(FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_willClear) begin
      FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_valueNext = 1'b0;
    end
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_1_write_mask = 1'b0;
    if(!when_MmuPlugin_l565) begin
      FetchL1Plugin_logic_translationStorage_logic_sl_1_write_mask = 1'b1;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
      end
      MmuPlugin_logic_refill_DONE_1 : begin
        FetchL1Plugin_logic_translationStorage_logic_sl_1_write_mask = (MmuPlugin_logic_refill_storageOhReg[0] ? 1'b1 : 1'b0);
        if(when_MmuPlugin_l505_2) begin
          FetchL1Plugin_logic_translationStorage_logic_sl_1_write_mask = 1'b0;
        end
      end
      MmuPlugin_logic_refill_DONE_2 : begin
        FetchL1Plugin_logic_translationStorage_logic_sl_1_write_mask = (MmuPlugin_logic_refill_storageOhReg[0] ? 1'b1 : 1'b0);
        if(when_MmuPlugin_l505_4) begin
          FetchL1Plugin_logic_translationStorage_logic_sl_1_write_mask = 1'b0;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_1_write_address = 5'bxxxxx;
    if(!when_MmuPlugin_l565) begin
      FetchL1Plugin_logic_translationStorage_logic_sl_1_write_address = MmuPlugin_logic_invalidate_counter;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
      end
      MmuPlugin_logic_refill_DONE_1 : begin
        FetchL1Plugin_logic_translationStorage_logic_sl_1_write_address = MmuPlugin_logic_refill_virtual[25 : 21];
      end
      MmuPlugin_logic_refill_DONE_2 : begin
        FetchL1Plugin_logic_translationStorage_logic_sl_1_write_address = MmuPlugin_logic_refill_virtual[25 : 21];
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_valid = 1'bx;
    if(!when_MmuPlugin_l565) begin
      FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_valid = 1'b0;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
      end
      MmuPlugin_logic_refill_DONE_1 : begin
        FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_valid = 1'b1;
      end
      MmuPlugin_logic_refill_DONE_2 : begin
        FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_valid = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_virtualAddress = 13'bxxxxxxxxxxxxx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
      end
      MmuPlugin_logic_refill_DONE_1 : begin
        FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_virtualAddress = MmuPlugin_logic_refill_virtual[38 : 26];
      end
      MmuPlugin_logic_refill_DONE_2 : begin
        FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_virtualAddress = MmuPlugin_logic_refill_virtual[38 : 26];
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_physicalAddress = 11'bxxxxxxxxxxx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
      end
      MmuPlugin_logic_refill_DONE_1 : begin
        FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_physicalAddress = _zz_FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_physicalAddress[10:0];
      end
      MmuPlugin_logic_refill_DONE_2 : begin
        FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_physicalAddress = _zz_FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_physicalAddress_1[10:0];
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowRead = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
      end
      MmuPlugin_logic_refill_DONE_1 : begin
        FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowRead = MmuPlugin_logic_refill_load_flags_R;
      end
      MmuPlugin_logic_refill_DONE_2 : begin
        FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowRead = MmuPlugin_logic_refill_load_flags_R;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowWrite = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
      end
      MmuPlugin_logic_refill_DONE_1 : begin
        FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowWrite = (MmuPlugin_logic_refill_load_flags_W && MmuPlugin_logic_refill_load_flags_D);
      end
      MmuPlugin_logic_refill_DONE_2 : begin
        FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowWrite = (MmuPlugin_logic_refill_load_flags_W && MmuPlugin_logic_refill_load_flags_D);
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowExecute = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
      end
      MmuPlugin_logic_refill_DONE_1 : begin
        FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowExecute = MmuPlugin_logic_refill_load_flags_X;
      end
      MmuPlugin_logic_refill_DONE_2 : begin
        FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowExecute = MmuPlugin_logic_refill_load_flags_X;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowUser = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
      end
      MmuPlugin_logic_refill_DONE_1 : begin
        FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowUser = MmuPlugin_logic_refill_load_flags_U;
      end
      MmuPlugin_logic_refill_DONE_2 : begin
        FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowUser = MmuPlugin_logic_refill_load_flags_U;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_1_allocId_willIncrement = 1'b0;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
      end
      MmuPlugin_logic_refill_DONE_1 : begin
        if(!when_MmuPlugin_l505_2) begin
          FetchL1Plugin_logic_translationStorage_logic_sl_1_allocId_willIncrement = 1'b1;
        end
      end
      MmuPlugin_logic_refill_DONE_2 : begin
        if(!when_MmuPlugin_l505_4) begin
          FetchL1Plugin_logic_translationStorage_logic_sl_1_allocId_willIncrement = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign FetchL1Plugin_logic_translationStorage_logic_sl_1_allocId_willClear = 1'b0;
  assign FetchL1Plugin_logic_translationStorage_logic_sl_1_allocId_willOverflowIfInc = 1'b1;
  assign FetchL1Plugin_logic_translationStorage_logic_sl_1_allocId_willOverflow = (FetchL1Plugin_logic_translationStorage_logic_sl_1_allocId_willOverflowIfInc && FetchL1Plugin_logic_translationStorage_logic_sl_1_allocId_willIncrement);
  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_0_write_mask = 3'b000;
    if(!when_MmuPlugin_l565) begin
      LsuPlugin_logic_translationStorage_logic_sl_0_write_mask = 3'b111;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
        LsuPlugin_logic_translationStorage_logic_sl_0_write_mask = _zz_LsuPlugin_logic_translationStorage_logic_sl_0_write_mask[2:0];
        if(when_MmuPlugin_l505_1) begin
          LsuPlugin_logic_translationStorage_logic_sl_0_write_mask = 3'b000;
        end
      end
      MmuPlugin_logic_refill_DONE_1 : begin
      end
      MmuPlugin_logic_refill_DONE_2 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_0_write_address = 5'bxxxxx;
    if(!when_MmuPlugin_l565) begin
      LsuPlugin_logic_translationStorage_logic_sl_0_write_address = MmuPlugin_logic_invalidate_counter;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
        LsuPlugin_logic_translationStorage_logic_sl_0_write_address = MmuPlugin_logic_refill_virtual[16 : 12];
      end
      MmuPlugin_logic_refill_DONE_1 : begin
      end
      MmuPlugin_logic_refill_DONE_2 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_0_write_data_valid = 1'bx;
    if(!when_MmuPlugin_l565) begin
      LsuPlugin_logic_translationStorage_logic_sl_0_write_data_valid = 1'b0;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
        LsuPlugin_logic_translationStorage_logic_sl_0_write_data_valid = 1'b1;
      end
      MmuPlugin_logic_refill_DONE_1 : begin
      end
      MmuPlugin_logic_refill_DONE_2 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_0_write_data_virtualAddress = 22'bxxxxxxxxxxxxxxxxxxxxxx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
        LsuPlugin_logic_translationStorage_logic_sl_0_write_data_virtualAddress = MmuPlugin_logic_refill_virtual[38 : 17];
      end
      MmuPlugin_logic_refill_DONE_1 : begin
      end
      MmuPlugin_logic_refill_DONE_2 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_0_write_data_physicalAddress = 20'bxxxxxxxxxxxxxxxxxxxx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
        LsuPlugin_logic_translationStorage_logic_sl_0_write_data_physicalAddress = _zz_LsuPlugin_logic_translationStorage_logic_sl_0_write_data_physicalAddress[19:0];
      end
      MmuPlugin_logic_refill_DONE_1 : begin
      end
      MmuPlugin_logic_refill_DONE_2 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowRead = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
        LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowRead = MmuPlugin_logic_refill_load_flags_R;
      end
      MmuPlugin_logic_refill_DONE_1 : begin
      end
      MmuPlugin_logic_refill_DONE_2 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowWrite = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
        LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowWrite = (MmuPlugin_logic_refill_load_flags_W && MmuPlugin_logic_refill_load_flags_D);
      end
      MmuPlugin_logic_refill_DONE_1 : begin
      end
      MmuPlugin_logic_refill_DONE_2 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowExecute = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
        LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowExecute = MmuPlugin_logic_refill_load_flags_X;
      end
      MmuPlugin_logic_refill_DONE_1 : begin
      end
      MmuPlugin_logic_refill_DONE_2 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowUser = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
        LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowUser = MmuPlugin_logic_refill_load_flags_U;
      end
      MmuPlugin_logic_refill_DONE_1 : begin
      end
      MmuPlugin_logic_refill_DONE_2 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_0_allocId_willIncrement = 1'b0;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
        if(!when_MmuPlugin_l505_1) begin
          LsuPlugin_logic_translationStorage_logic_sl_0_allocId_willIncrement = 1'b1;
        end
      end
      MmuPlugin_logic_refill_DONE_1 : begin
      end
      MmuPlugin_logic_refill_DONE_2 : begin
      end
      default : begin
      end
    endcase
  end

  assign LsuPlugin_logic_translationStorage_logic_sl_0_allocId_willClear = 1'b0;
  assign LsuPlugin_logic_translationStorage_logic_sl_0_allocId_willOverflowIfInc = (LsuPlugin_logic_translationStorage_logic_sl_0_allocId_value == 2'b10);
  assign LsuPlugin_logic_translationStorage_logic_sl_0_allocId_willOverflow = (LsuPlugin_logic_translationStorage_logic_sl_0_allocId_willOverflowIfInc && LsuPlugin_logic_translationStorage_logic_sl_0_allocId_willIncrement);
  always @(*) begin
    if(LsuPlugin_logic_translationStorage_logic_sl_0_allocId_willOverflow) begin
      LsuPlugin_logic_translationStorage_logic_sl_0_allocId_valueNext = 2'b00;
    end else begin
      LsuPlugin_logic_translationStorage_logic_sl_0_allocId_valueNext = (LsuPlugin_logic_translationStorage_logic_sl_0_allocId_value + _zz_LsuPlugin_logic_translationStorage_logic_sl_0_allocId_valueNext);
    end
    if(LsuPlugin_logic_translationStorage_logic_sl_0_allocId_willClear) begin
      LsuPlugin_logic_translationStorage_logic_sl_0_allocId_valueNext = 2'b00;
    end
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_1_write_mask = 1'b0;
    if(!when_MmuPlugin_l565) begin
      LsuPlugin_logic_translationStorage_logic_sl_1_write_mask = 1'b1;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
      end
      MmuPlugin_logic_refill_DONE_1 : begin
        LsuPlugin_logic_translationStorage_logic_sl_1_write_mask = (MmuPlugin_logic_refill_storageOhReg[1] ? 1'b1 : 1'b0);
        if(when_MmuPlugin_l505_3) begin
          LsuPlugin_logic_translationStorage_logic_sl_1_write_mask = 1'b0;
        end
      end
      MmuPlugin_logic_refill_DONE_2 : begin
        LsuPlugin_logic_translationStorage_logic_sl_1_write_mask = (MmuPlugin_logic_refill_storageOhReg[1] ? 1'b1 : 1'b0);
        if(when_MmuPlugin_l505_5) begin
          LsuPlugin_logic_translationStorage_logic_sl_1_write_mask = 1'b0;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_1_write_address = 5'bxxxxx;
    if(!when_MmuPlugin_l565) begin
      LsuPlugin_logic_translationStorage_logic_sl_1_write_address = MmuPlugin_logic_invalidate_counter;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
      end
      MmuPlugin_logic_refill_DONE_1 : begin
        LsuPlugin_logic_translationStorage_logic_sl_1_write_address = MmuPlugin_logic_refill_virtual[25 : 21];
      end
      MmuPlugin_logic_refill_DONE_2 : begin
        LsuPlugin_logic_translationStorage_logic_sl_1_write_address = MmuPlugin_logic_refill_virtual[25 : 21];
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_1_write_data_valid = 1'bx;
    if(!when_MmuPlugin_l565) begin
      LsuPlugin_logic_translationStorage_logic_sl_1_write_data_valid = 1'b0;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
      end
      MmuPlugin_logic_refill_DONE_1 : begin
        LsuPlugin_logic_translationStorage_logic_sl_1_write_data_valid = 1'b1;
      end
      MmuPlugin_logic_refill_DONE_2 : begin
        LsuPlugin_logic_translationStorage_logic_sl_1_write_data_valid = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_1_write_data_virtualAddress = 13'bxxxxxxxxxxxxx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
      end
      MmuPlugin_logic_refill_DONE_1 : begin
        LsuPlugin_logic_translationStorage_logic_sl_1_write_data_virtualAddress = MmuPlugin_logic_refill_virtual[38 : 26];
      end
      MmuPlugin_logic_refill_DONE_2 : begin
        LsuPlugin_logic_translationStorage_logic_sl_1_write_data_virtualAddress = MmuPlugin_logic_refill_virtual[38 : 26];
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_1_write_data_physicalAddress = 11'bxxxxxxxxxxx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
      end
      MmuPlugin_logic_refill_DONE_1 : begin
        LsuPlugin_logic_translationStorage_logic_sl_1_write_data_physicalAddress = _zz_LsuPlugin_logic_translationStorage_logic_sl_1_write_data_physicalAddress[10:0];
      end
      MmuPlugin_logic_refill_DONE_2 : begin
        LsuPlugin_logic_translationStorage_logic_sl_1_write_data_physicalAddress = _zz_LsuPlugin_logic_translationStorage_logic_sl_1_write_data_physicalAddress_1[10:0];
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowRead = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
      end
      MmuPlugin_logic_refill_DONE_1 : begin
        LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowRead = MmuPlugin_logic_refill_load_flags_R;
      end
      MmuPlugin_logic_refill_DONE_2 : begin
        LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowRead = MmuPlugin_logic_refill_load_flags_R;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowWrite = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
      end
      MmuPlugin_logic_refill_DONE_1 : begin
        LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowWrite = (MmuPlugin_logic_refill_load_flags_W && MmuPlugin_logic_refill_load_flags_D);
      end
      MmuPlugin_logic_refill_DONE_2 : begin
        LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowWrite = (MmuPlugin_logic_refill_load_flags_W && MmuPlugin_logic_refill_load_flags_D);
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowExecute = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
      end
      MmuPlugin_logic_refill_DONE_1 : begin
        LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowExecute = MmuPlugin_logic_refill_load_flags_X;
      end
      MmuPlugin_logic_refill_DONE_2 : begin
        LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowExecute = MmuPlugin_logic_refill_load_flags_X;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowUser = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
      end
      MmuPlugin_logic_refill_DONE_1 : begin
        LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowUser = MmuPlugin_logic_refill_load_flags_U;
      end
      MmuPlugin_logic_refill_DONE_2 : begin
        LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowUser = MmuPlugin_logic_refill_load_flags_U;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_1_allocId_willIncrement = 1'b0;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
      end
      MmuPlugin_logic_refill_DONE_1 : begin
        if(!when_MmuPlugin_l505_3) begin
          LsuPlugin_logic_translationStorage_logic_sl_1_allocId_willIncrement = 1'b1;
        end
      end
      MmuPlugin_logic_refill_DONE_2 : begin
        if(!when_MmuPlugin_l505_5) begin
          LsuPlugin_logic_translationStorage_logic_sl_1_allocId_willIncrement = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign LsuPlugin_logic_translationStorage_logic_sl_1_allocId_willClear = 1'b0;
  assign LsuPlugin_logic_translationStorage_logic_sl_1_allocId_willOverflowIfInc = 1'b1;
  assign LsuPlugin_logic_translationStorage_logic_sl_1_allocId_willOverflow = (LsuPlugin_logic_translationStorage_logic_sl_1_allocId_willOverflowIfInc && LsuPlugin_logic_translationStorage_logic_sl_1_allocId_willIncrement);
  assign MmuPlugin_logic_isMachine = (PrivilegedPlugin_logic_harts_0_privilege == 2'b11);
  assign MmuPlugin_logic_isSupervisor = (PrivilegedPlugin_logic_harts_0_privilege == 2'b01);
  assign MmuPlugin_logic_isUser = (PrivilegedPlugin_logic_harts_0_privilege == 2'b00);
  always @(*) begin
    MmuPlugin_api_fetchTranslationEnable = (MmuPlugin_logic_satp_mode == 4'b1000);
    if(MmuPlugin_logic_isMachine) begin
      MmuPlugin_api_fetchTranslationEnable = 1'b0;
    end
  end

  always @(*) begin
    MmuPlugin_api_lsuTranslationEnable = (MmuPlugin_logic_satp_mode == 4'b1000);
    if(when_MmuPlugin_l277) begin
      MmuPlugin_api_lsuTranslationEnable = 1'b0;
    end
    if(MmuPlugin_logic_isMachine) begin
      if(when_MmuPlugin_l279) begin
        MmuPlugin_api_lsuTranslationEnable = 1'b0;
      end
    end
  end

  assign when_MmuPlugin_l277 = ((! PrivilegedPlugin_logic_harts_0_m_status_mprv) && MmuPlugin_logic_isMachine);
  assign when_MmuPlugin_l279 = ((! PrivilegedPlugin_logic_harts_0_m_status_mprv) || (PrivilegedPlugin_logic_harts_0_m_status_mpp == 2'b11));
  assign LsuPlugin_logic_onAddress0_translationPort_logic_read_0_readAddress = execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0[16 : 12];
  assign _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_valid = LsuPlugin_logic_translationStorage_logic_sl_0_ways_0_spinal_port1;
  assign execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_valid = _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_valid[0];
  assign execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_virtualAddress = _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_valid[22 : 1];
  assign execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_physicalAddress = _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_valid[42 : 23];
  assign execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_allowRead = _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_valid[43];
  assign execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_allowWrite = _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_valid[44];
  assign execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_allowExecute = _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_valid[45];
  assign execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_allowUser = _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_valid[46];
  always @(*) begin
    execute_ctrl2_down_MMU_L0_HITS_PRE_VALID_lane0[0] = (execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_virtualAddress == execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0[38 : 17]);
    execute_ctrl2_down_MMU_L0_HITS_PRE_VALID_lane0[1] = (execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_virtualAddress == execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0[38 : 17]);
    execute_ctrl2_down_MMU_L0_HITS_PRE_VALID_lane0[2] = (execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_virtualAddress == execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0[38 : 17]);
  end

  always @(*) begin
    execute_ctrl3_down_MMU_L0_HITS_lane0[0] = (execute_ctrl3_down_MMU_L0_HITS_PRE_VALID_lane0[0] && execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_valid);
    execute_ctrl3_down_MMU_L0_HITS_lane0[1] = (execute_ctrl3_down_MMU_L0_HITS_PRE_VALID_lane0[1] && execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_valid);
    execute_ctrl3_down_MMU_L0_HITS_lane0[2] = (execute_ctrl3_down_MMU_L0_HITS_PRE_VALID_lane0[2] && execute_ctrl3_down_MMU_L0_ENTRIES_lane0_2_valid);
  end

  assign _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_valid = LsuPlugin_logic_translationStorage_logic_sl_0_ways_1_spinal_port1;
  assign execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_valid = _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_valid[0];
  assign execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_virtualAddress = _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_valid[22 : 1];
  assign execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_physicalAddress = _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_valid[42 : 23];
  assign execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_allowRead = _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_valid[43];
  assign execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_allowWrite = _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_valid[44];
  assign execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_allowExecute = _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_valid[45];
  assign execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_allowUser = _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_valid[46];
  assign _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_valid = LsuPlugin_logic_translationStorage_logic_sl_0_ways_2_spinal_port1;
  assign execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_valid = _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_valid[0];
  assign execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_virtualAddress = _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_valid[22 : 1];
  assign execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_physicalAddress = _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_valid[42 : 23];
  assign execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_allowRead = _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_valid[43];
  assign execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_allowWrite = _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_valid[44];
  assign execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_allowExecute = _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_valid[45];
  assign execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_allowUser = _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_valid[46];
  assign LsuPlugin_logic_onAddress0_translationPort_logic_read_1_readAddress = execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0[25 : 21];
  assign _zz_execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_valid = LsuPlugin_logic_translationStorage_logic_sl_1_ways_0_spinal_port1;
  assign execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_valid = _zz_execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_valid[0];
  assign execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_virtualAddress = _zz_execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_valid[13 : 1];
  assign execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_physicalAddress = _zz_execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_valid[24 : 14];
  assign execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_allowRead = _zz_execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_valid[25];
  assign execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_allowWrite = _zz_execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_valid[26];
  assign execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_allowExecute = _zz_execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_valid[27];
  assign execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_allowUser = _zz_execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_valid[28];
  assign execute_ctrl2_down_MMU_L1_HITS_PRE_VALID_lane0[0] = (execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_virtualAddress == execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0[38 : 26]);
  assign execute_ctrl3_down_MMU_L1_HITS_lane0[0] = (execute_ctrl3_down_MMU_L1_HITS_PRE_VALID_lane0[0] && execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_valid);
  assign LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits = {execute_ctrl3_down_MMU_L1_HITS_lane0,execute_ctrl3_down_MMU_L0_HITS_lane0};
  assign LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hit = (|LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits);
  assign _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_0 = LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits;
  assign LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_0 = _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_0[0];
  assign LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_1 = _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_0[1];
  assign LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_2 = _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_0[2];
  assign LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_3 = _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_0[3];
  always @(*) begin
    _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_oh[0] = (LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_0 && (! 1'b0));
    _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_oh[1] = (LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_1 && (! LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_0));
    _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_oh[2] = (LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_2 && (! LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_range_0_to_1));
    _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_oh[3] = (LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_3 && (! LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_range_0_to_2));
  end

  assign LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_range_0_to_1 = (|{LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_1,LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_0});
  assign LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_range_0_to_2 = (|{LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_2,{LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_1,LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_0}});
  assign LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_oh = _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_oh;
  assign _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute = LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_oh[0];
  assign _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_1 = LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_oh[1];
  assign _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_2 = LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_oh[2];
  assign _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_3 = LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_oh[3];
  assign LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute = _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_4[0];
  assign LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowRead = _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowRead[0];
  assign LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowWrite = _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowWrite[0];
  assign LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowUser = _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowUser[0];
  assign LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated = (((_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute ? {_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated,_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_1} : 32'h0) | (_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_1 ? {_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_2,_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_3} : 32'h0)) | ((_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_2 ? {_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_4,_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_5} : 32'h0) | (_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_3 ? {_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_6,_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_7} : 32'h0)));
  always @(*) begin
    LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_requireMmuLockup = MmuPlugin_api_lsuTranslationEnable;
    if(execute_ctrl3_down_LsuPlugin_logic_FORCE_PHYSICAL_lane0) begin
      LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_requireMmuLockup = 1'b0;
    end
  end

  always @(*) begin
    if(LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_requireMmuLockup) begin
      execute_ctrl3_down_MMU_HAZARD_lane0 = 1'b0;
    end else begin
      execute_ctrl3_down_MMU_HAZARD_lane0 = 1'b0;
    end
  end

  always @(*) begin
    if(LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_requireMmuLockup) begin
      execute_ctrl3_down_MMU_REFILL_lane0 = (! LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hit);
    end else begin
      execute_ctrl3_down_MMU_REFILL_lane0 = 1'b0;
    end
  end

  always @(*) begin
    if(LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_requireMmuLockup) begin
      execute_ctrl3_down_MMU_TRANSLATED_lane0 = LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated;
    end else begin
      execute_ctrl3_down_MMU_TRANSLATED_lane0 = execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[31:0];
    end
  end

  always @(*) begin
    if(LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_requireMmuLockup) begin
      execute_ctrl3_down_MMU_ALLOW_EXECUTE_lane0 = (LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute && (! (LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowUser && MmuPlugin_logic_isSupervisor)));
    end else begin
      execute_ctrl3_down_MMU_ALLOW_EXECUTE_lane0 = 1'b1;
    end
  end

  always @(*) begin
    if(LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_requireMmuLockup) begin
      execute_ctrl3_down_MMU_ALLOW_READ_lane0 = (LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowRead || (MmuPlugin_logic_status_mxr && LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute));
    end else begin
      execute_ctrl3_down_MMU_ALLOW_READ_lane0 = 1'b1;
    end
  end

  always @(*) begin
    if(LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_requireMmuLockup) begin
      execute_ctrl3_down_MMU_ALLOW_WRITE_lane0 = LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowWrite;
    end else begin
      execute_ctrl3_down_MMU_ALLOW_WRITE_lane0 = 1'b1;
    end
  end

  always @(*) begin
    if(LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_requireMmuLockup) begin
      execute_ctrl3_down_MMU_PAGE_FAULT_lane0 = (((LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowUser && MmuPlugin_logic_isSupervisor) && (! MmuPlugin_logic_status_sum)) || ((! LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowUser) && MmuPlugin_logic_isUser));
    end else begin
      execute_ctrl3_down_MMU_PAGE_FAULT_lane0 = 1'b0;
    end
  end

  always @(*) begin
    if(LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_requireMmuLockup) begin
      execute_ctrl3_down_MMU_ACCESS_FAULT_lane0 = 1'b0;
    end else begin
      execute_ctrl3_down_MMU_ACCESS_FAULT_lane0 = (execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[38 : 32] != 7'h0);
    end
  end

  assign execute_ctrl3_down_MMU_BYPASS_TRANSLATION_lane0 = (! LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_requireMmuLockup);
  assign execute_ctrl3_down_MMU_WAYS_OH_lane0 = LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_oh;
  assign execute_ctrl3_down_MMU_WAYS_PHYSICAL_lane0_0 = {execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_physicalAddress,execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[11 : 0]};
  assign execute_ctrl3_down_MMU_WAYS_PHYSICAL_lane0_1 = {execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_physicalAddress,execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[11 : 0]};
  assign execute_ctrl3_down_MMU_WAYS_PHYSICAL_lane0_2 = {execute_ctrl3_down_MMU_L0_ENTRIES_lane0_2_physicalAddress,execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[11 : 0]};
  assign execute_ctrl3_down_MMU_WAYS_PHYSICAL_lane0_3 = {execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_physicalAddress,execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[20 : 0]};
  assign FetchL1Plugin_logic_translationPort_logic_read_0_readAddress = fetch_logic_ctrls_1_down_Fetch_WORD_PC[16 : 12];
  assign _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_valid = FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_0_spinal_port1;
  assign fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_valid = _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_valid[0];
  assign fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_virtualAddress = _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_valid[22 : 1];
  assign fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_physicalAddress = _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_valid[42 : 23];
  assign fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_allowRead = _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_valid[43];
  assign fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_allowWrite = _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_valid[44];
  assign fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_allowExecute = _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_valid[45];
  assign fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_allowUser = _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_valid[46];
  always @(*) begin
    fetch_logic_ctrls_1_down_MMU_L0_HITS_PRE_VALID[0] = (fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_virtualAddress == fetch_logic_ctrls_1_down_Fetch_WORD_PC[38 : 17]);
    fetch_logic_ctrls_1_down_MMU_L0_HITS_PRE_VALID[1] = (fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_virtualAddress == fetch_logic_ctrls_1_down_Fetch_WORD_PC[38 : 17]);
  end

  always @(*) begin
    fetch_logic_ctrls_1_down_MMU_L0_HITS[0] = (fetch_logic_ctrls_1_down_MMU_L0_HITS_PRE_VALID[0] && fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_valid);
    fetch_logic_ctrls_1_down_MMU_L0_HITS[1] = (fetch_logic_ctrls_1_down_MMU_L0_HITS_PRE_VALID[1] && fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_valid);
  end

  assign _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_valid = FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_1_spinal_port1;
  assign fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_valid = _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_valid[0];
  assign fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_virtualAddress = _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_valid[22 : 1];
  assign fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_physicalAddress = _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_valid[42 : 23];
  assign fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_allowRead = _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_valid[43];
  assign fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_allowWrite = _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_valid[44];
  assign fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_allowExecute = _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_valid[45];
  assign fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_allowUser = _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_valid[46];
  assign FetchL1Plugin_logic_translationPort_logic_read_1_readAddress = fetch_logic_ctrls_1_down_Fetch_WORD_PC[25 : 21];
  assign _zz_fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_valid = FetchL1Plugin_logic_translationStorage_logic_sl_1_ways_0_spinal_port1;
  assign fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_valid = _zz_fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_valid[0];
  assign fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_virtualAddress = _zz_fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_valid[13 : 1];
  assign fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_physicalAddress = _zz_fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_valid[24 : 14];
  assign fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_allowRead = _zz_fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_valid[25];
  assign fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_allowWrite = _zz_fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_valid[26];
  assign fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_allowExecute = _zz_fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_valid[27];
  assign fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_allowUser = _zz_fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_valid[28];
  assign fetch_logic_ctrls_1_down_MMU_L1_HITS_PRE_VALID[0] = (fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_virtualAddress == fetch_logic_ctrls_1_down_Fetch_WORD_PC[38 : 26]);
  assign fetch_logic_ctrls_1_down_MMU_L1_HITS[0] = (fetch_logic_ctrls_1_down_MMU_L1_HITS_PRE_VALID[0] && fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_valid);
  assign FetchL1Plugin_logic_translationPort_logic_ctrl_hits = {fetch_logic_ctrls_1_down_MMU_L1_HITS,fetch_logic_ctrls_1_down_MMU_L0_HITS};
  assign FetchL1Plugin_logic_translationPort_logic_ctrl_hit = (|FetchL1Plugin_logic_translationPort_logic_ctrl_hits);
  assign _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_0 = FetchL1Plugin_logic_translationPort_logic_ctrl_hits;
  assign FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_0 = _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_0[0];
  assign FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_1 = _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_0[1];
  assign FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_2 = _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_0[2];
  always @(*) begin
    _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_oh[0] = (FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_0 && (! 1'b0));
    _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_oh[1] = (FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_1 && (! FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_0));
    _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_oh[2] = (FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_2 && (! FetchL1Plugin_logic_translationPort_logic_ctrl_hits_range_0_to_1));
  end

  assign FetchL1Plugin_logic_translationPort_logic_ctrl_hits_range_0_to_1 = (|{FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_1,FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_0});
  assign FetchL1Plugin_logic_translationPort_logic_ctrl_oh = _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_oh;
  assign _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute = FetchL1Plugin_logic_translationPort_logic_ctrl_oh[0];
  assign _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_1 = FetchL1Plugin_logic_translationPort_logic_ctrl_oh[1];
  assign _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_2 = FetchL1Plugin_logic_translationPort_logic_ctrl_oh[2];
  assign FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute = _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_3[0];
  assign FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowRead = _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowRead[0];
  assign FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowWrite = _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowWrite[0];
  assign FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowUser = _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowUser[0];
  assign FetchL1Plugin_logic_translationPort_logic_ctrl_lineTranslated = (((_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute ? {fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_physicalAddress,_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineTranslated} : 32'h0) | (_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_1 ? {fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_physicalAddress,_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineTranslated_1} : 32'h0)) | (_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_2 ? {fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_physicalAddress,fetch_logic_ctrls_1_down_Fetch_WORD_PC[20 : 0]} : 32'h0));
  always @(*) begin
    FetchL1Plugin_logic_translationPort_logic_ctrl_requireMmuLockup = MmuPlugin_api_fetchTranslationEnable;
    if(_zz_1) begin
      FetchL1Plugin_logic_translationPort_logic_ctrl_requireMmuLockup = 1'b0;
    end
  end

  always @(*) begin
    if(FetchL1Plugin_logic_translationPort_logic_ctrl_requireMmuLockup) begin
      fetch_logic_ctrls_1_down_MMU_HAZARD = 1'b0;
    end else begin
      fetch_logic_ctrls_1_down_MMU_HAZARD = 1'b0;
    end
  end

  always @(*) begin
    if(FetchL1Plugin_logic_translationPort_logic_ctrl_requireMmuLockup) begin
      fetch_logic_ctrls_1_down_MMU_REFILL = (! FetchL1Plugin_logic_translationPort_logic_ctrl_hit);
    end else begin
      fetch_logic_ctrls_1_down_MMU_REFILL = 1'b0;
    end
  end

  always @(*) begin
    if(FetchL1Plugin_logic_translationPort_logic_ctrl_requireMmuLockup) begin
      fetch_logic_ctrls_1_down_MMU_TRANSLATED = FetchL1Plugin_logic_translationPort_logic_ctrl_lineTranslated;
    end else begin
      fetch_logic_ctrls_1_down_MMU_TRANSLATED = fetch_logic_ctrls_1_down_Fetch_WORD_PC[31:0];
    end
  end

  always @(*) begin
    if(FetchL1Plugin_logic_translationPort_logic_ctrl_requireMmuLockup) begin
      fetch_logic_ctrls_1_down_MMU_ALLOW_EXECUTE = (FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute && (! (FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowUser && MmuPlugin_logic_isSupervisor)));
    end else begin
      fetch_logic_ctrls_1_down_MMU_ALLOW_EXECUTE = 1'b1;
    end
  end

  always @(*) begin
    if(FetchL1Plugin_logic_translationPort_logic_ctrl_requireMmuLockup) begin
      fetch_logic_ctrls_1_down_MMU_ALLOW_READ = (FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowRead || (MmuPlugin_logic_status_mxr && FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute));
    end else begin
      fetch_logic_ctrls_1_down_MMU_ALLOW_READ = 1'b1;
    end
  end

  always @(*) begin
    if(FetchL1Plugin_logic_translationPort_logic_ctrl_requireMmuLockup) begin
      fetch_logic_ctrls_1_down_MMU_ALLOW_WRITE = FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowWrite;
    end else begin
      fetch_logic_ctrls_1_down_MMU_ALLOW_WRITE = 1'b1;
    end
  end

  always @(*) begin
    if(FetchL1Plugin_logic_translationPort_logic_ctrl_requireMmuLockup) begin
      fetch_logic_ctrls_1_down_MMU_PAGE_FAULT = (((FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowUser && MmuPlugin_logic_isSupervisor) && (! MmuPlugin_logic_status_sum)) || ((! FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowUser) && MmuPlugin_logic_isUser));
    end else begin
      fetch_logic_ctrls_1_down_MMU_PAGE_FAULT = 1'b0;
    end
  end

  always @(*) begin
    if(FetchL1Plugin_logic_translationPort_logic_ctrl_requireMmuLockup) begin
      fetch_logic_ctrls_1_down_MMU_ACCESS_FAULT = 1'b0;
    end else begin
      fetch_logic_ctrls_1_down_MMU_ACCESS_FAULT = (fetch_logic_ctrls_1_down_Fetch_WORD_PC[38 : 32] != 7'h0);
    end
  end

  assign fetch_logic_ctrls_1_down_MMU_BYPASS_TRANSLATION = (! FetchL1Plugin_logic_translationPort_logic_ctrl_requireMmuLockup);
  assign fetch_logic_ctrls_1_down_MMU_WAYS_OH = FetchL1Plugin_logic_translationPort_logic_ctrl_oh;
  assign fetch_logic_ctrls_1_down_MMU_WAYS_PHYSICAL_0 = {fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_physicalAddress,fetch_logic_ctrls_1_down_Fetch_WORD_PC[11 : 0]};
  assign fetch_logic_ctrls_1_down_MMU_WAYS_PHYSICAL_1 = {fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_physicalAddress,fetch_logic_ctrls_1_down_Fetch_WORD_PC[11 : 0]};
  assign fetch_logic_ctrls_1_down_MMU_WAYS_PHYSICAL_2 = {fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_physicalAddress,fetch_logic_ctrls_1_down_Fetch_WORD_PC[20 : 0]};
  assign MmuPlugin_logic_refill_wantExit = 1'b0;
  always @(*) begin
    MmuPlugin_logic_refill_wantStart = 1'b0;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
      end
      MmuPlugin_logic_refill_DONE_1 : begin
      end
      MmuPlugin_logic_refill_DONE_2 : begin
      end
      default : begin
        MmuPlugin_logic_refill_wantStart = 1'b1;
      end
    endcase
  end

  assign MmuPlugin_logic_refill_wantKill = 1'b0;
  assign MmuPlugin_logic_refill_busy = (! (MmuPlugin_logic_refill_stateReg == MmuPlugin_logic_refill_IDLE));
  always @(*) begin
    MmuPlugin_logic_refill_cacheRefillAnySet = 1'b0;
    if(when_MmuPlugin_l400) begin
      MmuPlugin_logic_refill_cacheRefillAnySet = MmuPlugin_logic_accessBus_rsp_payload_waitAny;
    end
  end

  assign TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_cmd_ready = MmuPlugin_logic_refill_arbiter_io_inputs_0_ready;
  always @(*) begin
    MmuPlugin_logic_refill_arbiter_io_output_ready = 1'b0;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
        if(MmuPlugin_logic_refill_arbiter_io_output_valid) begin
          MmuPlugin_logic_refill_arbiter_io_output_ready = 1'b1;
        end
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
      end
      MmuPlugin_logic_refill_DONE_1 : begin
      end
      MmuPlugin_logic_refill_DONE_2 : begin
      end
      default : begin
      end
    endcase
  end

  assign MmuPlugin_logic_refill_events_onStorage_0_waiting = (MmuPlugin_logic_refill_busy && MmuPlugin_logic_refill_storageOhReg[0]);
  assign MmuPlugin_logic_refill_events_onStorage_1_waiting = (MmuPlugin_logic_refill_busy && MmuPlugin_logic_refill_storageOhReg[1]);
  assign MmuPlugin_logic_accessBus_rsp_toStream_valid = MmuPlugin_logic_accessBus_rsp_valid;
  assign MmuPlugin_logic_accessBus_rsp_toStream_payload_data = MmuPlugin_logic_accessBus_rsp_payload_data;
  assign MmuPlugin_logic_accessBus_rsp_toStream_payload_error = MmuPlugin_logic_accessBus_rsp_payload_error;
  assign MmuPlugin_logic_accessBus_rsp_toStream_payload_redo = MmuPlugin_logic_accessBus_rsp_payload_redo;
  assign MmuPlugin_logic_accessBus_rsp_toStream_payload_waitAny = MmuPlugin_logic_accessBus_rsp_payload_waitAny;
  always @(*) begin
    MmuPlugin_logic_accessBus_rsp_toStream_ready = MmuPlugin_logic_refill_load_rsp_ready;
    if(when_Stream_l477_2) begin
      MmuPlugin_logic_accessBus_rsp_toStream_ready = 1'b1;
    end
  end

  assign when_Stream_l477_2 = (! MmuPlugin_logic_refill_load_rsp_valid);
  assign MmuPlugin_logic_refill_load_rsp_valid = MmuPlugin_logic_accessBus_rsp_toStream_rValid;
  assign MmuPlugin_logic_refill_load_rsp_payload_data = MmuPlugin_logic_accessBus_rsp_toStream_rData_data;
  assign MmuPlugin_logic_refill_load_rsp_payload_error = MmuPlugin_logic_accessBus_rsp_toStream_rData_error;
  assign MmuPlugin_logic_refill_load_rsp_payload_redo = MmuPlugin_logic_accessBus_rsp_toStream_rData_redo;
  assign MmuPlugin_logic_refill_load_rsp_payload_waitAny = MmuPlugin_logic_accessBus_rsp_toStream_rData_waitAny;
  always @(*) begin
    MmuPlugin_logic_refill_load_rsp_ready = 1'b0;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            MmuPlugin_logic_refill_load_rsp_ready = 1'b1;
          end
        end
      end
      MmuPlugin_logic_refill_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            MmuPlugin_logic_refill_load_rsp_ready = 1'b1;
          end else begin
            if(!when_MmuPlugin_l534) begin
              MmuPlugin_logic_refill_load_rsp_ready = 1'b1;
            end
          end
        end
      end
      MmuPlugin_logic_refill_RSP_2 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            MmuPlugin_logic_refill_load_rsp_ready = 1'b1;
          end else begin
            if(!when_MmuPlugin_l534_1) begin
              MmuPlugin_logic_refill_load_rsp_ready = 1'b1;
            end
          end
        end
      end
      MmuPlugin_logic_refill_DONE_0 : begin
        MmuPlugin_logic_refill_load_rsp_ready = 1'b1;
      end
      MmuPlugin_logic_refill_DONE_1 : begin
        MmuPlugin_logic_refill_load_rsp_ready = 1'b1;
      end
      MmuPlugin_logic_refill_DONE_2 : begin
        MmuPlugin_logic_refill_load_rsp_ready = 1'b1;
      end
      default : begin
      end
    endcase
  end

  assign MmuPlugin_logic_refill_load_readed = MmuPlugin_logic_refill_load_rsp_payload_data[63 : 0];
  assign when_MmuPlugin_l400 = (MmuPlugin_logic_accessBus_rsp_valid && MmuPlugin_logic_accessBus_rsp_payload_redo);
  always @(*) begin
    MmuPlugin_logic_accessBus_cmd_valid = 1'b0;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
        if(when_MmuPlugin_l516) begin
          MmuPlugin_logic_accessBus_cmd_valid = 1'b1;
        end
      end
      MmuPlugin_logic_refill_CMD_1 : begin
        if(when_MmuPlugin_l516_1) begin
          MmuPlugin_logic_accessBus_cmd_valid = 1'b1;
        end
      end
      MmuPlugin_logic_refill_CMD_2 : begin
        if(when_MmuPlugin_l516_2) begin
          MmuPlugin_logic_accessBus_cmd_valid = 1'b1;
        end
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
      end
      MmuPlugin_logic_refill_DONE_1 : begin
      end
      MmuPlugin_logic_refill_DONE_2 : begin
      end
      default : begin
      end
    endcase
  end

  assign MmuPlugin_logic_accessBus_cmd_payload_address = MmuPlugin_logic_refill_load_address;
  assign MmuPlugin_logic_accessBus_cmd_payload_size = 2'b11;
  assign _zz_MmuPlugin_logic_refill_load_flags_V = MmuPlugin_logic_refill_load_readed;
  assign MmuPlugin_logic_refill_load_flags_V = _zz_MmuPlugin_logic_refill_load_flags_V[0];
  assign MmuPlugin_logic_refill_load_flags_R = _zz_MmuPlugin_logic_refill_load_flags_V[1];
  assign MmuPlugin_logic_refill_load_flags_W = _zz_MmuPlugin_logic_refill_load_flags_V[2];
  assign MmuPlugin_logic_refill_load_flags_X = _zz_MmuPlugin_logic_refill_load_flags_V[3];
  assign MmuPlugin_logic_refill_load_flags_U = _zz_MmuPlugin_logic_refill_load_flags_V[4];
  assign MmuPlugin_logic_refill_load_flags_G = _zz_MmuPlugin_logic_refill_load_flags_V[5];
  assign MmuPlugin_logic_refill_load_flags_A = _zz_MmuPlugin_logic_refill_load_flags_V[6];
  assign MmuPlugin_logic_refill_load_flags_D = _zz_MmuPlugin_logic_refill_load_flags_V[7];
  assign MmuPlugin_logic_refill_load_leaf = (MmuPlugin_logic_refill_load_flags_R || MmuPlugin_logic_refill_load_flags_X);
  assign MmuPlugin_logic_refill_load_reservedFault = (|(MmuPlugin_logic_refill_load_readed & 64'hffc0000000000000));
  always @(*) begin
    MmuPlugin_logic_refill_load_exception = (((((! MmuPlugin_logic_refill_load_flags_V) || ((! MmuPlugin_logic_refill_load_flags_R) && MmuPlugin_logic_refill_load_flags_W)) || MmuPlugin_logic_refill_load_rsp_payload_error) || ((! MmuPlugin_logic_refill_load_leaf) && ((MmuPlugin_logic_refill_load_flags_D || MmuPlugin_logic_refill_load_flags_A) || MmuPlugin_logic_refill_load_flags_U))) || MmuPlugin_logic_refill_load_reservedFault);
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
        if(when_MmuPlugin_l525) begin
          MmuPlugin_logic_refill_load_exception = 1'b1;
        end
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
      end
      MmuPlugin_logic_refill_DONE_1 : begin
      end
      MmuPlugin_logic_refill_DONE_2 : begin
      end
      default : begin
      end
    endcase
  end

  assign MmuPlugin_logic_refill_load_levelException_0 = 1'b0;
  always @(*) begin
    MmuPlugin_logic_refill_load_levelException_1 = 1'b0;
    if(when_MmuPlugin_l421) begin
      MmuPlugin_logic_refill_load_levelException_1 = 1'b1;
    end
  end

  always @(*) begin
    MmuPlugin_logic_refill_load_levelException_2 = 1'b0;
    if(when_MmuPlugin_l421_1) begin
      MmuPlugin_logic_refill_load_levelException_2 = 1'b1;
    end
    if(when_MmuPlugin_l421_2) begin
      MmuPlugin_logic_refill_load_levelException_2 = 1'b1;
    end
  end

  always @(*) begin
    MmuPlugin_logic_refill_load_nextLevelBase = 32'h0;
    MmuPlugin_logic_refill_load_nextLevelBase[20 : 12] = MmuPlugin_logic_refill_load_readed[18 : 10];
    MmuPlugin_logic_refill_load_nextLevelBase[29 : 21] = MmuPlugin_logic_refill_load_readed[27 : 19];
    MmuPlugin_logic_refill_load_nextLevelBase[31 : 30] = _zz_MmuPlugin_logic_refill_load_nextLevelBase[1:0];
  end

  always @(*) begin
    MmuPlugin_logic_refill_load_levelToPhysicalAddress_0 = 56'h0;
    MmuPlugin_logic_refill_load_levelToPhysicalAddress_0[20 : 12] = MmuPlugin_logic_refill_load_readed[18 : 10];
    MmuPlugin_logic_refill_load_levelToPhysicalAddress_0[29 : 21] = MmuPlugin_logic_refill_load_readed[27 : 19];
    MmuPlugin_logic_refill_load_levelToPhysicalAddress_0[55 : 30] = MmuPlugin_logic_refill_load_readed[53 : 28];
  end

  always @(*) begin
    MmuPlugin_logic_refill_load_levelToPhysicalAddress_1 = 56'h0;
    MmuPlugin_logic_refill_load_levelToPhysicalAddress_1[20 : 12] = MmuPlugin_logic_refill_virtual[20 : 12];
    MmuPlugin_logic_refill_load_levelToPhysicalAddress_1[29 : 21] = MmuPlugin_logic_refill_load_readed[27 : 19];
    MmuPlugin_logic_refill_load_levelToPhysicalAddress_1[55 : 30] = MmuPlugin_logic_refill_load_readed[53 : 28];
  end

  assign when_MmuPlugin_l421 = (MmuPlugin_logic_refill_load_readed[18 : 10] != 9'h0);
  always @(*) begin
    MmuPlugin_logic_refill_load_levelToPhysicalAddress_2 = 56'h0;
    MmuPlugin_logic_refill_load_levelToPhysicalAddress_2[20 : 12] = MmuPlugin_logic_refill_virtual[20 : 12];
    MmuPlugin_logic_refill_load_levelToPhysicalAddress_2[29 : 21] = MmuPlugin_logic_refill_virtual[29 : 21];
    MmuPlugin_logic_refill_load_levelToPhysicalAddress_2[55 : 30] = MmuPlugin_logic_refill_load_readed[53 : 28];
  end

  assign when_MmuPlugin_l421_1 = (MmuPlugin_logic_refill_load_readed[18 : 10] != 9'h0);
  assign when_MmuPlugin_l421_2 = (MmuPlugin_logic_refill_load_readed[27 : 19] != 9'h0);
  always @(*) begin
    TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_valid = 1'b0;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
        if(_zz_55) begin
          TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_valid = 1'b1;
        end
      end
      MmuPlugin_logic_refill_DONE_1 : begin
        if(_zz_55) begin
          TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_valid = 1'b1;
        end
      end
      MmuPlugin_logic_refill_DONE_2 : begin
        if(_zz_55) begin
          TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_valid = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    bits_pageFault = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
        bits_pageFault = MmuPlugin_logic_refill_fetch_0_pageFault;
      end
      MmuPlugin_logic_refill_DONE_1 : begin
        bits_pageFault = MmuPlugin_logic_refill_fetch_1_pageFault;
      end
      MmuPlugin_logic_refill_DONE_2 : begin
        bits_pageFault = MmuPlugin_logic_refill_fetch_2_pageFault;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    bits_accessFault = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
        bits_accessFault = MmuPlugin_logic_refill_fetch_0_accessFault;
      end
      MmuPlugin_logic_refill_DONE_1 : begin
        bits_accessFault = MmuPlugin_logic_refill_fetch_1_accessFault;
      end
      MmuPlugin_logic_refill_DONE_2 : begin
        bits_accessFault = MmuPlugin_logic_refill_fetch_2_accessFault;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    bits_pf = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
        bits_pf = MmuPlugin_logic_refill_fetch_0_pageFault;
      end
      MmuPlugin_logic_refill_DONE_1 : begin
        bits_pf = MmuPlugin_logic_refill_fetch_1_pageFault;
      end
      MmuPlugin_logic_refill_DONE_2 : begin
        bits_pf = MmuPlugin_logic_refill_fetch_2_pageFault;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    bits_ae_ptw = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
        bits_ae_ptw = (MmuPlugin_logic_refill_fetch_0_accessFault && (! MmuPlugin_logic_refill_load_leaf));
      end
      MmuPlugin_logic_refill_DONE_1 : begin
        bits_ae_ptw = (MmuPlugin_logic_refill_fetch_1_accessFault && (! MmuPlugin_logic_refill_load_leaf));
      end
      MmuPlugin_logic_refill_DONE_2 : begin
        bits_ae_ptw = (MmuPlugin_logic_refill_fetch_2_accessFault && (! MmuPlugin_logic_refill_load_leaf));
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    bits_ae_final = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
        bits_ae_final = (MmuPlugin_logic_refill_fetch_0_accessFault && MmuPlugin_logic_refill_load_leaf);
      end
      MmuPlugin_logic_refill_DONE_1 : begin
        bits_ae_final = (MmuPlugin_logic_refill_fetch_1_accessFault && MmuPlugin_logic_refill_load_leaf);
      end
      MmuPlugin_logic_refill_DONE_2 : begin
        bits_ae_final = (MmuPlugin_logic_refill_fetch_2_accessFault && MmuPlugin_logic_refill_load_leaf);
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    bits_level = 2'bxx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      MmuPlugin_logic_refill_RSP_2 : begin
      end
      MmuPlugin_logic_refill_DONE_0 : begin
        bits_level = 2'b10;
      end
      MmuPlugin_logic_refill_DONE_1 : begin
        bits_level = 2'b01;
      end
      MmuPlugin_logic_refill_DONE_2 : begin
        bits_level = 2'b00;
      end
      default : begin
      end
    endcase
  end

  assign bits_gf = 1'b0;
  assign bits_hr = 1'b0;
  assign bits_hw = 1'b0;
  assign bits_hx = 1'b0;
  assign bits_pte_d = MmuPlugin_logic_refill_load_flags_D;
  assign bits_pte_a = MmuPlugin_logic_refill_load_flags_A;
  assign bits_pte_g = MmuPlugin_logic_refill_load_flags_G;
  assign bits_pte_u = MmuPlugin_logic_refill_load_flags_U;
  assign bits_pte_x = MmuPlugin_logic_refill_load_flags_X;
  assign bits_pte_w = MmuPlugin_logic_refill_load_flags_W;
  assign bits_pte_r = MmuPlugin_logic_refill_load_flags_R;
  assign bits_pte_v = MmuPlugin_logic_refill_load_flags_V;
  assign bits_pte_ppn = _zz_bits_pte_ppn[19:0];
  assign MmuPlugin_logic_refill_fetch_0_pteFault = ((MmuPlugin_logic_refill_load_exception || MmuPlugin_logic_refill_load_levelException_0) || (! MmuPlugin_logic_refill_load_flags_A));
  assign MmuPlugin_logic_refill_fetch_0_leafAccessFault = (MmuPlugin_logic_refill_load_levelToPhysicalAddress_0[55 : 32] != 24'h0);
  assign MmuPlugin_logic_refill_fetch_0_pageFault = ((! MmuPlugin_logic_refill_load_rsp_payload_error) && MmuPlugin_logic_refill_fetch_0_pteFault);
  assign MmuPlugin_logic_refill_fetch_0_accessFault = (MmuPlugin_logic_refill_load_rsp_payload_error || ((! MmuPlugin_logic_refill_fetch_0_pteFault) && MmuPlugin_logic_refill_fetch_0_leafAccessFault));
  assign MmuPlugin_logic_refill_fetch_1_pteFault = ((MmuPlugin_logic_refill_load_exception || MmuPlugin_logic_refill_load_levelException_1) || (! MmuPlugin_logic_refill_load_flags_A));
  assign MmuPlugin_logic_refill_fetch_1_leafAccessFault = (MmuPlugin_logic_refill_load_levelToPhysicalAddress_1[55 : 32] != 24'h0);
  assign MmuPlugin_logic_refill_fetch_1_pageFault = ((! MmuPlugin_logic_refill_load_rsp_payload_error) && MmuPlugin_logic_refill_fetch_1_pteFault);
  assign MmuPlugin_logic_refill_fetch_1_accessFault = (MmuPlugin_logic_refill_load_rsp_payload_error || ((! MmuPlugin_logic_refill_fetch_1_pteFault) && MmuPlugin_logic_refill_fetch_1_leafAccessFault));
  assign MmuPlugin_logic_refill_fetch_2_pteFault = ((MmuPlugin_logic_refill_load_exception || MmuPlugin_logic_refill_load_levelException_2) || (! MmuPlugin_logic_refill_load_flags_A));
  assign MmuPlugin_logic_refill_fetch_2_leafAccessFault = (MmuPlugin_logic_refill_load_levelToPhysicalAddress_2[55 : 32] != 24'h0);
  assign MmuPlugin_logic_refill_fetch_2_pageFault = ((! MmuPlugin_logic_refill_load_rsp_payload_error) && MmuPlugin_logic_refill_fetch_2_pteFault);
  assign MmuPlugin_logic_refill_fetch_2_accessFault = (MmuPlugin_logic_refill_load_rsp_payload_error || ((! MmuPlugin_logic_refill_fetch_2_pteFault) && MmuPlugin_logic_refill_fetch_2_leafAccessFault));
  assign TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidate_cmd_ready = MmuPlugin_logic_invalidate_arbiter_io_inputs_0_ready;
  always @(*) begin
    MmuPlugin_logic_invalidate_arbiter_io_output_ready = 1'b0;
    if(!when_MmuPlugin_l565) begin
      if(when_MmuPlugin_l579) begin
        MmuPlugin_logic_invalidate_arbiter_io_output_ready = 1'b1;
      end
    end
  end

  assign when_MmuPlugin_l565 = (! MmuPlugin_logic_invalidate_busy);
  assign when_MmuPlugin_l579 = (&MmuPlugin_logic_invalidate_counter);
  always @(*) begin
    HistoryPlugin_logic_onFetch_valueNext = HistoryPlugin_logic_onFetch_value;
    if(HistoryPlugin_logic_onFetch_ports_0_valid) begin
      HistoryPlugin_logic_onFetch_valueNext = HistoryPlugin_logic_onFetch_ports_0_payload_history;
    end
    if(HistoryPlugin_logic_onFetch_ports_1_valid) begin
      HistoryPlugin_logic_onFetch_valueNext = HistoryPlugin_logic_onFetch_ports_1_payload_history;
    end
    if(HistoryPlugin_logic_onFetch_ports_2_valid) begin
      HistoryPlugin_logic_onFetch_valueNext = HistoryPlugin_logic_onFetch_ports_2_payload_history;
    end
  end

  assign HistoryPlugin_logic_onFetch_ports_0_valid = (|BtbPlugin_logic_historyPort_valid);
  assign HistoryPlugin_logic_onFetch_ports_0_payload_history = BtbPlugin_logic_historyPort_payload_history;
  assign HistoryPlugin_logic_onFetch_ports_1_valid = (|early0_BranchPlugin_logic_historyPort_valid);
  assign HistoryPlugin_logic_onFetch_ports_1_payload_history = early0_BranchPlugin_logic_historyPort_payload_history;
  assign HistoryPlugin_logic_onFetch_ports_2_valid = (|TrapPlugin_logic_harts_0_trap_historyPort_valid);
  assign HistoryPlugin_logic_onFetch_ports_2_payload_history = TrapPlugin_logic_harts_0_trap_historyPort_payload_history;
  assign fetch_logic_ctrls_0_down_Prediction_BRANCH_HISTORY = HistoryPlugin_logic_onFetch_valueNext;
  assign PerformanceCounterPlugin_logic_events_sums_0 = _zz_PerformanceCounterPlugin_logic_events_sums_0_1;
  assign PerformanceCounterPlugin_logic_events_sums_1 = _zz_PerformanceCounterPlugin_logic_events_sums_1_1;
  assign PerformanceCounterPlugin_logic_events_sums_2 = _zz_PerformanceCounterPlugin_logic_events_sums_2_1;
  assign PerformanceCounterPlugin_logic_events_sums_3 = _zz_PerformanceCounterPlugin_logic_events_sums_3_1;
  assign PerformanceCounterPlugin_logic_events_sums_4 = _zz_PerformanceCounterPlugin_logic_events_sums_4_1;
  assign PerformanceCounterPlugin_logic_events_sums_5 = _zz_PerformanceCounterPlugin_logic_events_sums_5_1;
  assign PerformanceCounterPlugin_logic_events_sums_6 = _zz_PerformanceCounterPlugin_logic_events_sums_6_1;
  assign PerformanceCounterPlugin_logic_events_sums_7 = _zz_PerformanceCounterPlugin_logic_events_sums_7_1;
  assign PerformanceCounterPlugin_logic_events_sums_8 = _zz_PerformanceCounterPlugin_logic_events_sums_8_1;
  assign PerformanceCounterPlugin_logic_events_sums_9 = _zz_PerformanceCounterPlugin_logic_events_sums_9_1;
  assign PerformanceCounterPlugin_logic_events_sums_10 = _zz_PerformanceCounterPlugin_logic_events_sums_10_1;
  assign PerformanceCounterPlugin_logic_events_sums_11 = _zz_PerformanceCounterPlugin_logic_events_sums_11_1;
  assign PerformanceCounterPlugin_logic_events_sums_12 = _zz_PerformanceCounterPlugin_logic_events_sums_12_1;
  assign PerformanceCounterPlugin_logic_events_sums_13 = _zz_PerformanceCounterPlugin_logic_events_sums_13_1;
  assign PerformanceCounterPlugin_logic_fsm_wantExit = 1'b0;
  always @(*) begin
    PerformanceCounterPlugin_logic_fsm_wantStart = 1'b0;
    case(PerformanceCounterPlugin_logic_fsm_stateReg)
      PerformanceCounterPlugin_logic_fsm_IDLE : begin
      end
      PerformanceCounterPlugin_logic_fsm_READ_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_CALC_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_CSR_WRITE : begin
      end
      default : begin
        PerformanceCounterPlugin_logic_fsm_wantStart = 1'b1;
      end
    endcase
  end

  assign PerformanceCounterPlugin_logic_fsm_wantKill = 1'b0;
  always @(*) begin
    PerformanceCounterPlugin_logic_fsm_csrReadCmd_ready = 1'b0;
    case(PerformanceCounterPlugin_logic_fsm_stateReg)
      PerformanceCounterPlugin_logic_fsm_IDLE : begin
        if(!PerformanceCounterPlugin_logic_fsm_csrWriteCmd_valid) begin
          if(!PerformanceCounterPlugin_logic_fsm_flusherCmd_valid) begin
            if(PerformanceCounterPlugin_logic_fsm_csrReadCmd_valid) begin
              PerformanceCounterPlugin_logic_fsm_csrReadCmd_ready = 1'b1;
            end
          end
        end
      end
      PerformanceCounterPlugin_logic_fsm_READ_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_CALC_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_CSR_WRITE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    PerformanceCounterPlugin_logic_fsm_flusherCmd_ready = 1'b0;
    case(PerformanceCounterPlugin_logic_fsm_stateReg)
      PerformanceCounterPlugin_logic_fsm_IDLE : begin
        if(!PerformanceCounterPlugin_logic_fsm_csrWriteCmd_valid) begin
          if(PerformanceCounterPlugin_logic_fsm_flusherCmd_valid) begin
            PerformanceCounterPlugin_logic_fsm_flusherCmd_ready = 1'b1;
          end
        end
      end
      PerformanceCounterPlugin_logic_fsm_READ_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_CALC_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_CSR_WRITE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    PerformanceCounterPlugin_logic_fsm_csrWriteCmd_ready = 1'b0;
    case(PerformanceCounterPlugin_logic_fsm_stateReg)
      PerformanceCounterPlugin_logic_fsm_IDLE : begin
      end
      PerformanceCounterPlugin_logic_fsm_READ_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_CALC_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_CSR_WRITE : begin
        PerformanceCounterPlugin_logic_fsm_csrWriteCmd_ready = 1'b1;
      end
      default : begin
      end
    endcase
  end

  assign _zz_PerformanceCounterPlugin_logic_fsm_cmd_address = PerformanceCounterPlugin_logic_fsm_cmd_oh[0];
  assign _zz_PerformanceCounterPlugin_logic_fsm_cmd_address_1 = PerformanceCounterPlugin_logic_fsm_cmd_oh[1];
  assign PerformanceCounterPlugin_logic_fsm_cmd_address = ((_zz_PerformanceCounterPlugin_logic_fsm_cmd_address ? 4'b0001 : 4'b0000) | (_zz_PerformanceCounterPlugin_logic_fsm_cmd_address_1 ? 4'b0000 : 4'b0000));
  always @(*) begin
    PerformanceCounterPlugin_logic_readPort_valid = 1'b0;
    case(PerformanceCounterPlugin_logic_fsm_stateReg)
      PerformanceCounterPlugin_logic_fsm_IDLE : begin
      end
      PerformanceCounterPlugin_logic_fsm_READ_LOW : begin
        PerformanceCounterPlugin_logic_readPort_valid = 1'b1;
      end
      PerformanceCounterPlugin_logic_fsm_CALC_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_CSR_WRITE : begin
      end
      default : begin
      end
    endcase
  end

  assign PerformanceCounterPlugin_logic_readPort_address = PerformanceCounterPlugin_logic_fsm_cmd_address;
  always @(*) begin
    PerformanceCounterPlugin_logic_writePort_valid = 1'b0;
    case(PerformanceCounterPlugin_logic_fsm_stateReg)
      PerformanceCounterPlugin_logic_fsm_IDLE : begin
      end
      PerformanceCounterPlugin_logic_fsm_READ_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_CALC_LOW : begin
        PerformanceCounterPlugin_logic_writePort_valid = 1'b1;
      end
      PerformanceCounterPlugin_logic_fsm_CSR_WRITE : begin
      end
      default : begin
      end
    endcase
  end

  assign PerformanceCounterPlugin_logic_writePort_address = PerformanceCounterPlugin_logic_readPort_address;
  always @(*) begin
    PerformanceCounterPlugin_logic_writePort_data = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(PerformanceCounterPlugin_logic_fsm_stateReg)
      PerformanceCounterPlugin_logic_fsm_IDLE : begin
      end
      PerformanceCounterPlugin_logic_fsm_READ_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_CALC_LOW : begin
        PerformanceCounterPlugin_logic_writePort_data = _zz_PerformanceCounterPlugin_logic_writePort_data[63:0];
      end
      PerformanceCounterPlugin_logic_fsm_CSR_WRITE : begin
      end
      default : begin
      end
    endcase
  end

  assign PerformanceCounterPlugin_logic_fsm_calc_a = {PerformanceCounterPlugin_logic_fsm_ramReaded[63 : 7],_zz_PerformanceCounterPlugin_logic_fsm_calc_a};
  assign PerformanceCounterPlugin_logic_fsm_calc_b = ({7'd0,PerformanceCounterPlugin_logic_fsm_counterReaded[7]} <<< 3'd7);
  assign PerformanceCounterPlugin_logic_fsm_calc_sum = ({1'b0,PerformanceCounterPlugin_logic_fsm_calc_a} + _zz_PerformanceCounterPlugin_logic_fsm_calc_sum);
  assign PerformanceCounterPlugin_logic_fsm_idleCsrAddress = (PerformanceCounterPlugin_logic_fsm_csrReadCmd_valid ? PerformanceCounterPlugin_logic_fsm_csrReadCmd_payload_address : PerformanceCounterPlugin_logic_fsm_csrWriteCmd_payload_address);
  always @(*) begin
    PerformanceCounterPlugin_logic_fsm_holdCsrWrite = 1'b1;
    case(PerformanceCounterPlugin_logic_fsm_stateReg)
      PerformanceCounterPlugin_logic_fsm_IDLE : begin
        PerformanceCounterPlugin_logic_fsm_holdCsrWrite = 1'b0;
      end
      PerformanceCounterPlugin_logic_fsm_READ_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_CALC_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_CSR_WRITE : begin
        PerformanceCounterPlugin_logic_fsm_holdCsrWrite = 1'b0;
      end
      default : begin
      end
    endcase
  end

  assign PerformanceCounterPlugin_logic_flusher_hits = {PerformanceCounterPlugin_logic_counters_instret_needFlush,PerformanceCounterPlugin_logic_counters_cycle_needFlush};
  assign PerformanceCounterPlugin_logic_flusher_hit = (|PerformanceCounterPlugin_logic_flusher_hits);
  assign PerformanceCounterPlugin_logic_flusher_hits_ohFirst_input = PerformanceCounterPlugin_logic_flusher_hits;
  assign PerformanceCounterPlugin_logic_flusher_hits_ohFirst_masked = (PerformanceCounterPlugin_logic_flusher_hits_ohFirst_input & (~ _zz_PerformanceCounterPlugin_logic_flusher_hits_ohFirst_masked));
  assign PerformanceCounterPlugin_logic_flusher_oh = PerformanceCounterPlugin_logic_flusher_hits_ohFirst_masked;
  assign PerformanceCounterPlugin_logic_fsm_flusherCmd_valid = PerformanceCounterPlugin_logic_flusher_hit;
  assign PerformanceCounterPlugin_logic_fsm_flusherCmd_payload_oh = PerformanceCounterPlugin_logic_flusher_oh;
  assign PerformanceCounterPlugin_logic_csrDecode_addr = CsrAccessPlugin_bus_decode_address[1 : 0];
  always @(*) begin
    PerformanceCounterPlugin_logic_csrDecode_mok = 1'bx;
    case(PerformanceCounterPlugin_logic_csrDecode_addr)
      2'b00 : begin
        PerformanceCounterPlugin_logic_csrDecode_mok = PerformanceCounterPlugin_logic_counters_cycle_mcounteren;
      end
      2'b10 : begin
        PerformanceCounterPlugin_logic_csrDecode_mok = PerformanceCounterPlugin_logic_counters_instret_mcounteren;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    PerformanceCounterPlugin_logic_csrDecode_sok = 1'bx;
    case(PerformanceCounterPlugin_logic_csrDecode_addr)
      2'b00 : begin
        PerformanceCounterPlugin_logic_csrDecode_sok = PerformanceCounterPlugin_logic_counters_cycle_scounteren;
      end
      2'b10 : begin
        PerformanceCounterPlugin_logic_csrDecode_sok = PerformanceCounterPlugin_logic_counters_instret_scounteren;
      end
      default : begin
      end
    endcase
  end

  assign PerformanceCounterPlugin_logic_csrDecode_privOk = (&(PrivilegedPlugin_logic_harts_0_privilege | {PerformanceCounterPlugin_logic_csrDecode_mok,PerformanceCounterPlugin_logic_csrDecode_sok}));
  assign PerformanceCounterPlugin_logic_fsm_csrReadCmd_fire = (PerformanceCounterPlugin_logic_fsm_csrReadCmd_valid && PerformanceCounterPlugin_logic_fsm_csrReadCmd_ready);
  assign PerformanceCounterPlugin_logic_csrRead_requested = (CsrAccessPlugin_bus_read_valid && REG_CSR_PerformanceCounterPlugin_logic_csrFilter);
  assign PerformanceCounterPlugin_logic_fsm_csrReadCmd_valid = (PerformanceCounterPlugin_logic_csrRead_requested && (! PerformanceCounterPlugin_logic_csrRead_fired));
  assign PerformanceCounterPlugin_logic_fsm_csrReadCmd_payload_address = CsrAccessPlugin_bus_read_address[1 : 0];
  assign when_PerformanceCounterPlugin_l342 = ((! PerformanceCounterPlugin_logic_csrRead_fired) || (! PerformanceCounterPlugin_logic_fsm_done));
  assign PerformanceCounterPlugin_logic_fsm_csrWriteCmd_fire = (PerformanceCounterPlugin_logic_fsm_csrWriteCmd_valid && PerformanceCounterPlugin_logic_fsm_csrWriteCmd_ready);
  always @(*) begin
    PerformanceCounterPlugin_logic_fsm_csrWriteCmd_valid = 1'b0;
    if(when_CsrAccessPlugin_l349_3) begin
      if(when_PerformanceCounterPlugin_l357) begin
        PerformanceCounterPlugin_logic_fsm_csrWriteCmd_valid = 1'b1;
      end
    end
  end

  assign PerformanceCounterPlugin_logic_fsm_csrWriteCmd_payload_address = CsrAccessPlugin_bus_write_address[1 : 0];
  assign fetch_logic_flushes_0_doIt = (|{(DecoderPlugin_logic_laneLogic_0_flushPort_valid && 1'b1),{(early0_EnvPlugin_logic_flushPort_valid && 1'b1),{(CsrAccessPlugin_logic_flushPort_valid && 1'b1),{(early0_BranchPlugin_logic_flushPort_valid && 1'b1),{(LsuPlugin_logic_flushPort_valid && 1'b1),((BtbPlugin_logic_flushPort_valid && _zz_fetch_logic_flushes_0_doIt) && (_zz_fetch_logic_flushes_0_doIt_1 || _zz_fetch_logic_flushes_0_doIt_2))}}}}});
  assign fetch_logic_ctrls_1_throwWhen_FetchPipelinePlugin_l48 = fetch_logic_flushes_0_doIt;
  assign fetch_logic_flushes_1_doIt = (|{(DecoderPlugin_logic_laneLogic_0_flushPort_valid && 1'b1),{(early0_EnvPlugin_logic_flushPort_valid && 1'b1),{(CsrAccessPlugin_logic_flushPort_valid && 1'b1),{(early0_BranchPlugin_logic_flushPort_valid && 1'b1),(LsuPlugin_logic_flushPort_valid && 1'b1)}}}});
  assign fetch_logic_ctrls_2_forgetsSingleRequest_FetchPipelinePlugin_l50 = fetch_logic_flushes_1_doIt;
  assign CsrAccessPlugin_logic_fsm_wantExit = 1'b0;
  always @(*) begin
    CsrAccessPlugin_logic_fsm_wantStart = 1'b0;
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_READ : begin
      end
      CsrAccessPlugin_logic_fsm_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_COMPLETION : begin
      end
      default : begin
        CsrAccessPlugin_logic_fsm_wantStart = 1'b1;
      end
    endcase
  end

  assign CsrAccessPlugin_logic_fsm_wantKill = 1'b0;
  always @(*) begin
    CsrAccessPlugin_logic_fsm_interface_fire = 1'b0;
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_READ : begin
      end
      CsrAccessPlugin_logic_fsm_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_COMPLETION : begin
        if(execute_ctrl2_down_isReady) begin
          CsrAccessPlugin_logic_fsm_interface_fire = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign CsrAccessPlugin_logic_fsm_inject_csrAddress = execute_ctrl2_down_Decode_UOP_lane0[31 : 20];
  assign CsrAccessPlugin_logic_fsm_inject_immZero = (execute_ctrl2_down_Decode_UOP_lane0[19 : 15] == 5'h0);
  assign CsrAccessPlugin_logic_fsm_inject_srcZero = (execute_ctrl2_down_CsrAccessPlugin_CSR_IMM_lane0 ? CsrAccessPlugin_logic_fsm_inject_immZero : (execute_ctrl2_down_Decode_UOP_lane0[19 : 15] == 5'h0));
  assign CsrAccessPlugin_logic_fsm_inject_csrWrite = (! (execute_ctrl2_down_CsrAccessPlugin_CSR_MASK_lane0 && CsrAccessPlugin_logic_fsm_inject_srcZero));
  assign CsrAccessPlugin_logic_fsm_inject_csrRead = (! ((! execute_ctrl2_down_CsrAccessPlugin_CSR_MASK_lane0) && (! execute_ctrl2_up_RD_ENABLE_lane0)));
  assign COMB_CSR_768 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h300);
  assign COMB_CSR_256 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h100);
  assign COMB_CSR_384 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h180);
  assign COMB_CSR_944 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h3b0);
  assign COMB_CSR_928 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h3a0);
  assign COMB_CSR_945 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h3b1);
  assign COMB_CSR_946 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h3b2);
  assign COMB_CSR_947 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h3b3);
  assign COMB_CSR_PmpPlugin_logic_allFilter = (|{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h3a2),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h3a0),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h3bf),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h3be),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == _zz_COMB_CSR_PmpPlugin_logic_allFilter),{_zz_COMB_CSR_PmpPlugin_logic_allFilter_1,{_zz_COMB_CSR_PmpPlugin_logic_allFilter_2,_zz_COMB_CSR_PmpPlugin_logic_allFilter_3}}}}}}});
  assign COMB_CSR_794 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h31a);
  assign COMB_CSR_1952 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h7a0);
  assign COMB_CSR_1953 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h7a1);
  assign COMB_CSR_1954 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h7a2);
  assign COMB_CSR_3857 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hf11);
  assign COMB_CSR_3858 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hf12);
  assign COMB_CSR_3859 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hf13);
  assign COMB_CSR_3860 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hf14);
  assign COMB_CSR_769 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h301);
  assign COMB_CSR_834 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h342);
  assign COMB_CSR_836 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h344);
  assign COMB_CSR_772 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h304);
  assign COMB_CSR_770 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h302);
  assign COMB_CSR_771 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h303);
  assign COMB_CSR_4016 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hfb0);
  assign COMB_CSR_774 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h306);
  assign COMB_CSR_322 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h142);
  assign COMB_CSR_778 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h30a);
  assign COMB_CSR_260 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h104);
  assign COMB_CSR_324 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h144);
  assign COMB_CSR_3504 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hdb0);
  assign COMB_CSR_3073 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc01);
  assign COMB_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_tvecFilter = (|{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h105),(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h305)});
  assign COMB_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_epcFilter = (|{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h141),(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h341)});
  assign COMB_CSR_262 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h106);
  assign COMB_CSR_800 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h320);
  assign COMB_CSR_UNAMED_1 = (|{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h33f),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc1f),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb1f),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h33e),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc1e),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb1e),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == _zz_COMB_CSR_UNAMED_1),{_zz_COMB_CSR_UNAMED_1_1,{_zz_COMB_CSR_UNAMED_1_2,_zz_COMB_CSR_UNAMED_1_3}}}}}}}}});
  assign COMB_CSR_266 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h10a);
  assign COMB_CSR_CsrRamPlugin_csrMapper_selFilter = (|{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc02),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb02),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc00),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb00),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h140),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h141),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == _zz_COMB_CSR_CsrRamPlugin_csrMapper_selFilter),{_zz_COMB_CSR_CsrRamPlugin_csrMapper_selFilter_1,{_zz_COMB_CSR_CsrRamPlugin_csrMapper_selFilter_2,_zz_COMB_CSR_CsrRamPlugin_csrMapper_selFilter_3}}}}}}}}});
  assign COMB_CSR_PerformanceCounterPlugin_logic_csrFilter = (|{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc02),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb02),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc00),(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb00)}}});
  assign COMB_CSR_CsrAccessPlugin_logic_trapNextOnWriteFilter = (|{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h100),(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h300)});
  assign CsrAccessPlugin_logic_fsm_inject_implemented = (|{COMB_CSR_CsrAccessPlugin_logic_trapNextOnWriteFilter,{COMB_CSR_PerformanceCounterPlugin_logic_csrFilter,{COMB_CSR_CsrRamPlugin_csrMapper_selFilter,{COMB_CSR_266,{COMB_CSR_UNAMED_1,{COMB_CSR_800,{COMB_CSR_262,{COMB_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_epcFilter,{COMB_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_tvecFilter,{COMB_CSR_3073,{_zz_CsrAccessPlugin_logic_fsm_inject_implemented,_zz_CsrAccessPlugin_logic_fsm_inject_implemented_1}}}}}}}}}}});
  assign CsrAccessPlugin_logic_fsm_inject_onDecodeDo = ((execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_down_CsrAccessPlugin_SEL_lane0) && (CsrAccessPlugin_logic_fsm_stateReg == CsrAccessPlugin_logic_fsm_IDLE));
  assign when_CsrAccessPlugin_l157 = (CsrAccessPlugin_logic_fsm_inject_onDecodeDo && COMB_CSR_384);
  assign when_MmuPlugin_l223 = (PrivilegedPlugin_logic_harts_0_m_status_tvm && (PrivilegedPlugin_logic_harts_0_privilege == 2'b01));
  assign when_CsrAccessPlugin_l157_1 = (CsrAccessPlugin_logic_fsm_inject_onDecodeDo && COMB_CSR_PmpPlugin_logic_allFilter);
  assign when_CsrAccessPlugin_l157_2 = (CsrAccessPlugin_logic_fsm_inject_onDecodeDo && COMB_CSR_794);
  assign when_CsrService_l121 = (! 1'b1);
  assign when_CsrAccessPlugin_l157_3 = (CsrAccessPlugin_logic_fsm_inject_onDecodeDo && COMB_CSR_1952);
  assign when_CsrService_l121_1 = (! 1'b1);
  assign when_CsrAccessPlugin_l157_4 = (CsrAccessPlugin_logic_fsm_inject_onDecodeDo && COMB_CSR_1953);
  assign when_CsrService_l121_2 = (! 1'b1);
  assign when_CsrAccessPlugin_l157_5 = (CsrAccessPlugin_logic_fsm_inject_onDecodeDo && COMB_CSR_1954);
  assign when_CsrService_l121_3 = (! 1'b1);
  assign when_CsrAccessPlugin_l157_6 = (CsrAccessPlugin_logic_fsm_inject_onDecodeDo && COMB_CSR_3073);
  assign when_CsrService_l198 = (when_CsrService_l232 || when_CsrService_l210);
  assign when_CsrService_l199 = (! PrivilegedPlugin_logic_harts_0_time_accessable);
  assign when_CsrAccessPlugin_l157_7 = (CsrAccessPlugin_logic_fsm_inject_onDecodeDo && COMB_CSR_UNAMED_1);
  assign when_CsrService_l121_4 = (! 1'b1);
  assign when_CsrAccessPlugin_l157_8 = (CsrAccessPlugin_logic_fsm_inject_onDecodeDo && COMB_CSR_CsrRamPlugin_csrMapper_selFilter);
  assign when_CsrService_l121_5 = (! 1'b1);
  assign when_CsrAccessPlugin_l157_9 = (CsrAccessPlugin_logic_fsm_inject_onDecodeDo && COMB_CSR_PerformanceCounterPlugin_logic_csrFilter);
  assign when_PerformanceCounterPlugin_l327 = (CsrAccessPlugin_bus_decode_address[9 : 8] == 2'b00);
  assign when_PerformanceCounterPlugin_l328 = (CsrAccessPlugin_bus_decode_write || (! PerformanceCounterPlugin_logic_csrDecode_privOk));
  assign when_CsrAccessPlugin_l157_10 = (CsrAccessPlugin_logic_fsm_inject_onDecodeDo && COMB_CSR_CsrAccessPlugin_logic_trapNextOnWriteFilter);
  assign CsrAccessPlugin_logic_fsm_inject_trap = ((! CsrAccessPlugin_logic_fsm_inject_implemented) || CsrAccessPlugin_bus_decode_exception);
  assign CsrAccessPlugin_bus_decode_read = CsrAccessPlugin_logic_fsm_inject_csrRead;
  assign CsrAccessPlugin_bus_decode_write = CsrAccessPlugin_logic_fsm_inject_csrWrite;
  assign CsrAccessPlugin_bus_decode_address = CsrAccessPlugin_logic_fsm_inject_csrAddress;
  assign CsrAccessPlugin_logic_fsm_interface_uopId = execute_ctrl2_down_Decode_UOP_ID_lane0;
  assign CsrAccessPlugin_logic_fsm_interface_rs1 = execute_ctrl2_up_integer_RS1_lane0;
  assign CsrAccessPlugin_logic_fsm_interface_uop = execute_ctrl2_down_Decode_UOP_lane0;
  assign CsrAccessPlugin_logic_fsm_interface_doImm = execute_ctrl2_down_CsrAccessPlugin_CSR_IMM_lane0;
  assign CsrAccessPlugin_logic_fsm_interface_doMask = execute_ctrl2_down_CsrAccessPlugin_CSR_MASK_lane0;
  assign CsrAccessPlugin_logic_fsm_interface_doClear = execute_ctrl2_down_CsrAccessPlugin_CSR_CLEAR_lane0;
  assign CsrAccessPlugin_logic_fsm_interface_rdEnable = execute_ctrl2_up_RD_ENABLE_lane0;
  assign CsrAccessPlugin_logic_fsm_interface_rdPhys = execute_ctrl2_down_RD_PHYS_lane0;
  assign CsrAccessPlugin_logic_fsm_inject_freeze = ((execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_down_CsrAccessPlugin_SEL_lane0) && (! CsrAccessPlugin_logic_fsm_inject_unfreeze));
  always @(*) begin
    CsrAccessPlugin_logic_flushPort_valid = 1'b0;
    if(CsrAccessPlugin_logic_fsm_inject_flushReg) begin
      CsrAccessPlugin_logic_flushPort_valid = 1'b1;
    end
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_READ : begin
      end
      CsrAccessPlugin_logic_fsm_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_COMPLETION : begin
      end
      default : begin
        if(CsrAccessPlugin_logic_fsm_inject_onDecodeDo) begin
          if(CsrAccessPlugin_logic_fsm_inject_sampled) begin
            if(CsrAccessPlugin_logic_fsm_inject_trapReg) begin
              CsrAccessPlugin_logic_flushPort_valid = 1'b1;
            end else begin
              if(CsrAccessPlugin_logic_fsm_inject_busTrapReg) begin
                CsrAccessPlugin_logic_flushPort_valid = 1'b1;
              end
            end
          end
        end
      end
    endcase
  end

  assign CsrAccessPlugin_logic_flushPort_payload_uopId = execute_ctrl2_down_Decode_UOP_ID_lane0;
  assign CsrAccessPlugin_logic_flushPort_payload_self = 1'b0;
  always @(*) begin
    CsrAccessPlugin_logic_trapPort_valid = 1'b0;
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_READ : begin
      end
      CsrAccessPlugin_logic_fsm_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_COMPLETION : begin
      end
      default : begin
        if(CsrAccessPlugin_logic_fsm_inject_onDecodeDo) begin
          if(CsrAccessPlugin_logic_fsm_inject_sampled) begin
            if(CsrAccessPlugin_logic_fsm_inject_trapReg) begin
              CsrAccessPlugin_logic_trapPort_valid = 1'b1;
            end else begin
              if(CsrAccessPlugin_logic_fsm_inject_busTrapReg) begin
                CsrAccessPlugin_logic_trapPort_valid = 1'b1;
              end
            end
          end
        end
      end
    endcase
  end

  always @(*) begin
    CsrAccessPlugin_logic_trapPort_payload_exception = 1'b1;
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_READ : begin
      end
      CsrAccessPlugin_logic_fsm_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_COMPLETION : begin
      end
      default : begin
        if(CsrAccessPlugin_logic_fsm_inject_onDecodeDo) begin
          if(CsrAccessPlugin_logic_fsm_inject_sampled) begin
            if(!CsrAccessPlugin_logic_fsm_inject_trapReg) begin
              if(CsrAccessPlugin_logic_fsm_inject_busTrapReg) begin
                CsrAccessPlugin_logic_trapPort_payload_exception = 1'b0;
              end
            end
          end
        end
      end
    endcase
  end

  always @(*) begin
    CsrAccessPlugin_logic_trapPort_payload_code = 4'b0010;
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_READ : begin
      end
      CsrAccessPlugin_logic_fsm_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_COMPLETION : begin
      end
      default : begin
        if(CsrAccessPlugin_logic_fsm_inject_onDecodeDo) begin
          if(CsrAccessPlugin_logic_fsm_inject_sampled) begin
            if(!CsrAccessPlugin_logic_fsm_inject_trapReg) begin
              if(CsrAccessPlugin_logic_fsm_inject_busTrapReg) begin
                CsrAccessPlugin_logic_trapPort_payload_code = CsrAccessPlugin_logic_fsm_inject_busTrapCodeReg;
              end
            end
          end
        end
      end
    endcase
  end

  assign CsrAccessPlugin_logic_trapPort_payload_tval = {7'd0, execute_ctrl2_down_Decode_UOP_lane0};
  assign CsrAccessPlugin_logic_trapPort_payload_arg = 3'b000;
  assign when_CsrAccessPlugin_l199 = (! execute_freeze_valid);
  always @(*) begin
    CsrAccessPlugin_logic_fsm_readLogic_onReadsDo = 1'b0;
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_READ : begin
        CsrAccessPlugin_logic_fsm_readLogic_onReadsDo = CsrAccessPlugin_logic_fsm_interface_read;
      end
      CsrAccessPlugin_logic_fsm_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_COMPLETION : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    CsrAccessPlugin_logic_fsm_readLogic_onReadsFireDo = 1'b0;
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_READ : begin
        if(when_CsrAccessPlugin_l302) begin
          CsrAccessPlugin_logic_fsm_readLogic_onReadsFireDo = CsrAccessPlugin_logic_fsm_interface_read;
        end
      end
      CsrAccessPlugin_logic_fsm_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_COMPLETION : begin
      end
      default : begin
      end
    endcase
  end

  assign CsrAccessPlugin_bus_read_valid = CsrAccessPlugin_logic_fsm_readLogic_onReadsDo;
  assign CsrAccessPlugin_bus_read_address = CsrAccessPlugin_logic_fsm_interface_uop[31 : 20];
  assign CsrAccessPlugin_bus_read_moving = (! CsrAccessPlugin_bus_read_halt);
  assign when_CsrAccessPlugin_l258 = (CsrAccessPlugin_logic_fsm_readLogic_onReadsDo && REG_CSR_CsrRamPlugin_csrMapper_selFilter);
  assign CsrAccessPlugin_logic_fsm_readLogic_csrValue = (((((_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_32 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_43) | (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_53 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_64)) | ((_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_75 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_86) | (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_97 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_108))) | (((_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_119 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_128) | (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_133 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_143)) | ((_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_154 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_164) | (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_175 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_186)))) | ((((_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_197 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_208) | (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_219 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_228)) | ((_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_239 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_249) | (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_260 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_271))) | (((_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_282 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_291) | (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_302 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_313)) | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_322)));
  assign CsrAccessPlugin_bus_read_data = CsrAccessPlugin_logic_fsm_readLogic_csrValue;
  always @(*) begin
    CsrAccessPlugin_bus_read_toWriteBits = CsrAccessPlugin_logic_fsm_readLogic_csrValue;
    if(when_CsrAccessPlugin_l285) begin
      if(when_CsrService_l232) begin
        CsrAccessPlugin_bus_read_toWriteBits[9 : 9] = PrivilegedPlugin_logic_harts_0_s_ip_seipSoft;
      end
    end
  end

  assign when_CsrAccessPlugin_l285 = (CsrAccessPlugin_logic_fsm_readLogic_onReadsDo && REG_CSR_836);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue = REG_CSR_768;
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_1 = REG_CSR_256;
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_2 = REG_CSR_384;
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3 = REG_CSR_944;
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5 = REG_CSR_928;
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_6 = REG_CSR_945;
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_8 = REG_CSR_946;
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_10 = REG_CSR_947;
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_14 = REG_CSR_836;
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_16 = REG_CSR_772;
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_19 = REG_CSR_771;
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_22 = REG_CSR_774;
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_25 = REG_CSR_778;
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_29 = REG_CSR_262;
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_30 = REG_CSR_800;
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_31 = REG_CSR_266;
  assign when_CsrService_l232 = 1'b1;
  assign CsrAccessPlugin_bus_write_moving = (! CsrAccessPlugin_bus_write_halt);
  assign CsrAccessPlugin_logic_fsm_writeLogic_alu_mask = (CsrAccessPlugin_logic_fsm_interface_doImm ? _zz_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask : CsrAccessPlugin_logic_fsm_interface_rs1);
  assign CsrAccessPlugin_logic_fsm_writeLogic_alu_masked = (CsrAccessPlugin_logic_fsm_interface_doClear ? (CsrAccessPlugin_logic_fsm_interface_aluInput & (~ CsrAccessPlugin_logic_fsm_writeLogic_alu_mask)) : (CsrAccessPlugin_logic_fsm_interface_aluInput | CsrAccessPlugin_logic_fsm_writeLogic_alu_mask));
  assign CsrAccessPlugin_logic_fsm_writeLogic_alu_result = (CsrAccessPlugin_logic_fsm_interface_doMask ? CsrAccessPlugin_logic_fsm_writeLogic_alu_masked : CsrAccessPlugin_logic_fsm_writeLogic_alu_mask);
  always @(*) begin
    CsrAccessPlugin_bus_write_bits = CsrAccessPlugin_logic_fsm_writeLogic_alu_result;
    if(when_CsrAccessPlugin_l349) begin
      CsrAccessPlugin_bus_write_bits[1 : 0] = 2'b00;
    end
    if(when_CsrAccessPlugin_l349_1) begin
      CsrAccessPlugin_bus_write_bits[0 : 0] = 1'b0;
    end
  end

  assign CsrAccessPlugin_bus_write_address = CsrAccessPlugin_logic_fsm_interface_uop[31 : 20];
  always @(*) begin
    CsrAccessPlugin_logic_fsm_writeLogic_onWritesDo = 1'b0;
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_READ : begin
      end
      CsrAccessPlugin_logic_fsm_WRITE : begin
        CsrAccessPlugin_logic_fsm_writeLogic_onWritesDo = CsrAccessPlugin_logic_fsm_interface_write;
      end
      CsrAccessPlugin_logic_fsm_COMPLETION : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo = 1'b0;
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_READ : begin
      end
      CsrAccessPlugin_logic_fsm_WRITE : begin
        if(when_CsrAccessPlugin_l331) begin
          CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo = CsrAccessPlugin_logic_fsm_interface_write;
        end
      end
      CsrAccessPlugin_logic_fsm_COMPLETION : begin
      end
      default : begin
      end
    endcase
  end

  assign CsrAccessPlugin_bus_write_valid = CsrAccessPlugin_logic_fsm_writeLogic_onWritesDo;
  assign when_CsrService_l210 = 1'b1;
  assign when_CsrAccessPlugin_l352 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_768);
  assign switch_PrivilegedPlugin_l581 = CsrAccessPlugin_bus_write_bits[12 : 11];
  assign when_CsrAccessPlugin_l352_1 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_256);
  assign when_CsrAccessPlugin_l359 = ((|((MmuPlugin_logic_satpModeWrite != 4'b0000) && (MmuPlugin_logic_satpModeWrite != 4'b1000))) == 1'b0);
  assign when_CsrAccessPlugin_l352_2 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_384);
  assign when_CsrAccessPlugin_l359_1 = ((|PmpPlugin_logic_entries_0_isLocked) == 1'b0);
  assign when_CsrAccessPlugin_l352_3 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_944);
  assign when_CsrAccessPlugin_l352_4 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_928);
  assign when_CsrAccessPlugin_l359_2 = ((|PmpPlugin_logic_entries_1_isLocked) == 1'b0);
  assign when_CsrAccessPlugin_l352_5 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_945);
  assign when_CsrAccessPlugin_l359_3 = ((|PmpPlugin_logic_entries_2_isLocked) == 1'b0);
  assign when_CsrAccessPlugin_l352_6 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_946);
  assign when_CsrAccessPlugin_l359_4 = ((|PmpPlugin_logic_entries_3_isLocked) == 1'b0);
  assign when_CsrAccessPlugin_l352_7 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_947);
  assign when_CsrAccessPlugin_l352_8 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_834);
  assign when_CsrAccessPlugin_l352_9 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_836);
  assign when_CsrAccessPlugin_l352_10 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_772);
  assign when_CsrAccessPlugin_l352_11 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_770);
  assign when_CsrAccessPlugin_l352_12 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_771);
  assign when_CsrAccessPlugin_l352_13 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_774);
  assign when_CsrAccessPlugin_l352_14 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_322);
  assign when_CsrAccessPlugin_l352_15 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_778);
  assign when_CsrAccessPlugin_l352_16 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_260);
  assign when_CsrAccessPlugin_l352_17 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_324);
  assign when_CsrAccessPlugin_l349 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesDo && REG_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_tvecFilter);
  assign when_CsrAccessPlugin_l349_1 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesDo && REG_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_epcFilter);
  assign when_CsrAccessPlugin_l352_18 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_262);
  assign when_CsrAccessPlugin_l352_19 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_800);
  assign when_CsrAccessPlugin_l352_20 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_266);
  assign when_CsrAccessPlugin_l349_2 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesDo && REG_CSR_CsrRamPlugin_csrMapper_selFilter);
  assign when_CsrAccessPlugin_l349_3 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesDo && REG_CSR_PerformanceCounterPlugin_logic_csrFilter);
  assign when_PerformanceCounterPlugin_l357 = (! PerformanceCounterPlugin_logic_csrWrite_fired);
  assign when_PerformanceCounterPlugin_l359 = (! PerformanceCounterPlugin_logic_fsm_csrWriteCmd_ready);
  assign CsrAccessPlugin_logic_wbWi_valid = execute_ctrl3_down_CsrAccessPlugin_SEL_lane0;
  assign CsrAccessPlugin_logic_wbWi_payload = CsrAccessPlugin_logic_fsm_interface_csrValue;
  assign CsrRamPlugin_logic_writeLogic_hits = {CsrRamPlugin_setup_initPort_valid,{CsrRamPlugin_csrMapper_write_valid,{TrapPlugin_logic_harts_0_crsPorts_write_valid,PerformanceCounterPlugin_logic_writePort_valid}}};
  assign CsrRamPlugin_logic_writeLogic_hit = (|CsrRamPlugin_logic_writeLogic_hits);
  assign CsrRamPlugin_logic_writeLogic_hits_ohFirst_input = CsrRamPlugin_logic_writeLogic_hits;
  assign CsrRamPlugin_logic_writeLogic_hits_ohFirst_masked = (CsrRamPlugin_logic_writeLogic_hits_ohFirst_input & (~ _zz_CsrRamPlugin_logic_writeLogic_hits_ohFirst_masked));
  assign CsrRamPlugin_logic_writeLogic_oh = CsrRamPlugin_logic_writeLogic_hits_ohFirst_masked;
  assign _zz_PerformanceCounterPlugin_logic_writePort_ready = CsrRamPlugin_logic_writeLogic_oh[0];
  assign _zz_TrapPlugin_logic_harts_0_crsPorts_write_ready = CsrRamPlugin_logic_writeLogic_oh[1];
  assign _zz_CsrRamPlugin_csrMapper_write_ready = CsrRamPlugin_logic_writeLogic_oh[2];
  assign _zz_CsrRamPlugin_setup_initPort_ready = CsrRamPlugin_logic_writeLogic_oh[3];
  assign CsrRamPlugin_logic_writeLogic_port_valid = CsrRamPlugin_logic_writeLogic_hit;
  assign CsrRamPlugin_logic_writeLogic_port_payload_address = (((_zz_PerformanceCounterPlugin_logic_writePort_ready ? PerformanceCounterPlugin_logic_writePort_address : 4'b0000) | (_zz_TrapPlugin_logic_harts_0_crsPorts_write_ready ? TrapPlugin_logic_harts_0_crsPorts_write_address : 4'b0000)) | ((_zz_CsrRamPlugin_csrMapper_write_ready ? CsrRamPlugin_csrMapper_write_address : 4'b0000) | (_zz_CsrRamPlugin_setup_initPort_ready ? CsrRamPlugin_setup_initPort_address : 4'b0000)));
  assign CsrRamPlugin_logic_writeLogic_port_payload_data = (((_zz_PerformanceCounterPlugin_logic_writePort_ready ? PerformanceCounterPlugin_logic_writePort_data : 64'h0) | (_zz_TrapPlugin_logic_harts_0_crsPorts_write_ready ? TrapPlugin_logic_harts_0_crsPorts_write_data : 64'h0)) | ((_zz_CsrRamPlugin_csrMapper_write_ready ? CsrRamPlugin_csrMapper_write_data : 64'h0) | (_zz_CsrRamPlugin_setup_initPort_ready ? CsrRamPlugin_setup_initPort_data : 64'h0)));
  assign PerformanceCounterPlugin_logic_writePort_ready = _zz_PerformanceCounterPlugin_logic_writePort_ready;
  assign TrapPlugin_logic_harts_0_crsPorts_write_ready = _zz_TrapPlugin_logic_harts_0_crsPorts_write_ready;
  assign CsrRamPlugin_csrMapper_write_ready = _zz_CsrRamPlugin_csrMapper_write_ready;
  assign CsrRamPlugin_setup_initPort_ready = _zz_CsrRamPlugin_setup_initPort_ready;
  assign CsrRamPlugin_logic_readLogic_hits = {CsrRamPlugin_csrMapper_read_valid,{TrapPlugin_logic_harts_0_crsPorts_read_valid,PerformanceCounterPlugin_logic_readPort_valid}};
  assign CsrRamPlugin_logic_readLogic_hit = (|CsrRamPlugin_logic_readLogic_hits);
  assign CsrRamPlugin_logic_readLogic_hits_ohFirst_input = CsrRamPlugin_logic_readLogic_hits;
  assign CsrRamPlugin_logic_readLogic_hits_ohFirst_masked = (CsrRamPlugin_logic_readLogic_hits_ohFirst_input & (~ _zz_CsrRamPlugin_logic_readLogic_hits_ohFirst_masked));
  assign CsrRamPlugin_logic_readLogic_oh = CsrRamPlugin_logic_readLogic_hits_ohFirst_masked;
  assign _zz_CsrRamPlugin_logic_readLogic_sel = CsrRamPlugin_logic_readLogic_oh[1];
  assign _zz_CsrRamPlugin_logic_readLogic_sel_1 = CsrRamPlugin_logic_readLogic_oh[2];
  assign CsrRamPlugin_logic_readLogic_sel = {_zz_CsrRamPlugin_logic_readLogic_sel_1,_zz_CsrRamPlugin_logic_readLogic_sel};
  assign CsrRamPlugin_logic_readLogic_port_rsp = CsrRamPlugin_logic_mem_spinal_port1;
  assign CsrRamPlugin_logic_readLogic_port_cmd_valid = (((|CsrRamPlugin_logic_readLogic_oh) && (! CsrRamPlugin_logic_writeLogic_port_valid)) && (! CsrRamPlugin_logic_readLogic_busy));
  assign CsrRamPlugin_logic_readLogic_port_cmd_payload = _zz_CsrRamPlugin_logic_readLogic_port_cmd_payload;
  assign PerformanceCounterPlugin_logic_readPort_ready = CsrRamPlugin_logic_readLogic_ohReg[0];
  assign TrapPlugin_logic_harts_0_crsPorts_read_ready = CsrRamPlugin_logic_readLogic_ohReg[1];
  assign CsrRamPlugin_csrMapper_read_ready = CsrRamPlugin_logic_readLogic_ohReg[2];
  assign PerformanceCounterPlugin_logic_readPort_data = CsrRamPlugin_logic_readLogic_port_rsp;
  assign TrapPlugin_logic_harts_0_crsPorts_read_data = CsrRamPlugin_logic_readLogic_port_rsp;
  assign CsrRamPlugin_csrMapper_read_data = CsrRamPlugin_logic_readLogic_port_rsp;
  assign CsrRamPlugin_logic_flush_done = CsrRamPlugin_logic_flush_counter[4];
  assign CsrRamPlugin_setup_initPort_valid = (! CsrRamPlugin_logic_flush_done);
  assign CsrRamPlugin_setup_initPort_address = CsrRamPlugin_logic_flush_counter[3:0];
  assign CsrRamPlugin_setup_initPort_data = 64'h0;
  assign execute_lane0_bypasser_integer_RS1_port_valid = (! execute_freeze_valid);
  assign execute_lane0_bypasser_integer_RS1_port_address = execute_ctrl0_down_RS1_PHYS_lane0[4 : 0];
  always @(*) begin
    execute_lane0_bypasser_integer_RS1_bypassEnables[0] = (((execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_up_RD_ENABLE_lane0) && (execute_ctrl2_down_RD_PHYS_lane0 == execute_ctrl1_down_RS1_PHYS_lane0)) && 1'b1);
    execute_lane0_bypasser_integer_RS1_bypassEnables[1] = (((execute_ctrl3_up_LANE_SEL_lane0 && execute_ctrl3_up_RD_ENABLE_lane0) && (execute_ctrl3_down_RD_PHYS_lane0 == execute_ctrl1_down_RS1_PHYS_lane0)) && 1'b1);
    execute_lane0_bypasser_integer_RS1_bypassEnables[2] = (((execute_ctrl4_up_LANE_SEL_lane0 && execute_ctrl4_up_RD_ENABLE_lane0) && (execute_ctrl4_down_RD_PHYS_lane0 == execute_ctrl1_down_RS1_PHYS_lane0)) && 1'b1);
    execute_lane0_bypasser_integer_RS1_bypassEnables[3] = (((execute_ctrl5_up_LANE_SEL_lane0 && execute_ctrl5_up_RD_ENABLE_lane0) && (execute_ctrl5_down_RD_PHYS_lane0 == execute_ctrl1_down_RS1_PHYS_lane0)) && 1'b1);
    execute_lane0_bypasser_integer_RS1_bypassEnables[4] = 1'b1;
  end

  assign _zz_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0 = execute_lane0_bypasser_integer_RS1_bypassEnables;
  assign execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0 = _zz_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0[0];
  assign execute_lane0_bypasser_integer_RS1_bypassEnables_bools_1 = _zz_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0[1];
  assign execute_lane0_bypasser_integer_RS1_bypassEnables_bools_2 = _zz_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0[2];
  assign execute_lane0_bypasser_integer_RS1_bypassEnables_bools_3 = _zz_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0[3];
  assign execute_lane0_bypasser_integer_RS1_bypassEnables_bools_4 = _zz_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0[4];
  always @(*) begin
    _zz_execute_lane0_bypasser_integer_RS1_sel[0] = (execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0 && (! 1'b0));
    _zz_execute_lane0_bypasser_integer_RS1_sel[1] = (execute_lane0_bypasser_integer_RS1_bypassEnables_bools_1 && (! execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0));
    _zz_execute_lane0_bypasser_integer_RS1_sel[2] = (execute_lane0_bypasser_integer_RS1_bypassEnables_bools_2 && (! execute_lane0_bypasser_integer_RS1_bypassEnables_range_0_to_1));
    _zz_execute_lane0_bypasser_integer_RS1_sel[3] = (execute_lane0_bypasser_integer_RS1_bypassEnables_bools_3 && (! execute_lane0_bypasser_integer_RS1_bypassEnables_range_0_to_2));
    _zz_execute_lane0_bypasser_integer_RS1_sel[4] = (execute_lane0_bypasser_integer_RS1_bypassEnables_bools_4 && (! execute_lane0_bypasser_integer_RS1_bypassEnables_range_0_to_3));
  end

  assign execute_lane0_bypasser_integer_RS1_bypassEnables_range_0_to_1 = (|{execute_lane0_bypasser_integer_RS1_bypassEnables_bools_1,execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0});
  assign execute_lane0_bypasser_integer_RS1_bypassEnables_range_0_to_2 = (|{execute_lane0_bypasser_integer_RS1_bypassEnables_bools_2,{execute_lane0_bypasser_integer_RS1_bypassEnables_bools_1,execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0}});
  assign execute_lane0_bypasser_integer_RS1_bypassEnables_range_0_to_3 = (|{execute_lane0_bypasser_integer_RS1_bypassEnables_bools_3,{execute_lane0_bypasser_integer_RS1_bypassEnables_bools_2,{execute_lane0_bypasser_integer_RS1_bypassEnables_bools_1,execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0}}});
  assign execute_lane0_bypasser_integer_RS1_sel = _zz_execute_lane0_bypasser_integer_RS1_sel;
  assign _zz_execute_ctrl1_down_integer_RS1_lane0 = execute_lane0_bypasser_integer_RS1_sel[4 : 1];
  always @(*) begin
    _zz_execute_ctrl1_down_integer_RS1_lane0_1 = (((_zz_execute_ctrl1_down_integer_RS1_lane0[0] ? execute_ctrl3_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : 64'h0) | (_zz_execute_ctrl1_down_integer_RS1_lane0[1] ? execute_ctrl4_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : 64'h0)) | ((_zz_execute_ctrl1_down_integer_RS1_lane0[2] ? execute_ctrl5_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : 64'h0) | (_zz_execute_ctrl1_down_integer_RS1_lane0[3] ? execute_lane0_bypasser_integer_RS1_port_data : 64'h0)));
    if(when_ExecuteLanePlugin_l196) begin
      _zz_execute_ctrl1_down_integer_RS1_lane0_1 = execute_ctrl2_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
    end
  end

  assign execute_ctrl1_down_integer_RS1_lane0 = _zz_execute_ctrl1_down_integer_RS1_lane0_1;
  assign when_ExecuteLanePlugin_l196 = execute_lane0_bypasser_integer_RS1_sel[0];
  assign execute_lane0_bypasser_integer_RS2_port_valid = (! execute_freeze_valid);
  assign execute_lane0_bypasser_integer_RS2_port_address = execute_ctrl0_down_RS2_PHYS_lane0[4 : 0];
  always @(*) begin
    execute_lane0_bypasser_integer_RS2_bypassEnables[0] = (((execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_up_RD_ENABLE_lane0) && (execute_ctrl2_down_RD_PHYS_lane0 == execute_ctrl1_down_RS2_PHYS_lane0)) && 1'b1);
    execute_lane0_bypasser_integer_RS2_bypassEnables[1] = (((execute_ctrl3_up_LANE_SEL_lane0 && execute_ctrl3_up_RD_ENABLE_lane0) && (execute_ctrl3_down_RD_PHYS_lane0 == execute_ctrl1_down_RS2_PHYS_lane0)) && 1'b1);
    execute_lane0_bypasser_integer_RS2_bypassEnables[2] = (((execute_ctrl4_up_LANE_SEL_lane0 && execute_ctrl4_up_RD_ENABLE_lane0) && (execute_ctrl4_down_RD_PHYS_lane0 == execute_ctrl1_down_RS2_PHYS_lane0)) && 1'b1);
    execute_lane0_bypasser_integer_RS2_bypassEnables[3] = (((execute_ctrl5_up_LANE_SEL_lane0 && execute_ctrl5_up_RD_ENABLE_lane0) && (execute_ctrl5_down_RD_PHYS_lane0 == execute_ctrl1_down_RS2_PHYS_lane0)) && 1'b1);
    execute_lane0_bypasser_integer_RS2_bypassEnables[4] = 1'b1;
  end

  assign _zz_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0 = execute_lane0_bypasser_integer_RS2_bypassEnables;
  assign execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0 = _zz_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0[0];
  assign execute_lane0_bypasser_integer_RS2_bypassEnables_bools_1 = _zz_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0[1];
  assign execute_lane0_bypasser_integer_RS2_bypassEnables_bools_2 = _zz_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0[2];
  assign execute_lane0_bypasser_integer_RS2_bypassEnables_bools_3 = _zz_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0[3];
  assign execute_lane0_bypasser_integer_RS2_bypassEnables_bools_4 = _zz_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0[4];
  always @(*) begin
    _zz_execute_lane0_bypasser_integer_RS2_sel[0] = (execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0 && (! 1'b0));
    _zz_execute_lane0_bypasser_integer_RS2_sel[1] = (execute_lane0_bypasser_integer_RS2_bypassEnables_bools_1 && (! execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0));
    _zz_execute_lane0_bypasser_integer_RS2_sel[2] = (execute_lane0_bypasser_integer_RS2_bypassEnables_bools_2 && (! execute_lane0_bypasser_integer_RS2_bypassEnables_range_0_to_1));
    _zz_execute_lane0_bypasser_integer_RS2_sel[3] = (execute_lane0_bypasser_integer_RS2_bypassEnables_bools_3 && (! execute_lane0_bypasser_integer_RS2_bypassEnables_range_0_to_2));
    _zz_execute_lane0_bypasser_integer_RS2_sel[4] = (execute_lane0_bypasser_integer_RS2_bypassEnables_bools_4 && (! execute_lane0_bypasser_integer_RS2_bypassEnables_range_0_to_3));
  end

  assign execute_lane0_bypasser_integer_RS2_bypassEnables_range_0_to_1 = (|{execute_lane0_bypasser_integer_RS2_bypassEnables_bools_1,execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0});
  assign execute_lane0_bypasser_integer_RS2_bypassEnables_range_0_to_2 = (|{execute_lane0_bypasser_integer_RS2_bypassEnables_bools_2,{execute_lane0_bypasser_integer_RS2_bypassEnables_bools_1,execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0}});
  assign execute_lane0_bypasser_integer_RS2_bypassEnables_range_0_to_3 = (|{execute_lane0_bypasser_integer_RS2_bypassEnables_bools_3,{execute_lane0_bypasser_integer_RS2_bypassEnables_bools_2,{execute_lane0_bypasser_integer_RS2_bypassEnables_bools_1,execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0}}});
  assign execute_lane0_bypasser_integer_RS2_sel = _zz_execute_lane0_bypasser_integer_RS2_sel;
  assign _zz_execute_ctrl1_down_integer_RS2_lane0 = execute_lane0_bypasser_integer_RS2_sel[4 : 1];
  always @(*) begin
    _zz_execute_ctrl1_down_integer_RS2_lane0_1 = (((_zz_execute_ctrl1_down_integer_RS2_lane0[0] ? execute_ctrl3_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : 64'h0) | (_zz_execute_ctrl1_down_integer_RS2_lane0[1] ? execute_ctrl4_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : 64'h0)) | ((_zz_execute_ctrl1_down_integer_RS2_lane0[2] ? execute_ctrl5_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : 64'h0) | (_zz_execute_ctrl1_down_integer_RS2_lane0[3] ? execute_lane0_bypasser_integer_RS2_port_data : 64'h0)));
    if(when_ExecuteLanePlugin_l196_1) begin
      _zz_execute_ctrl1_down_integer_RS2_lane0_1 = execute_ctrl2_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
    end
  end

  assign execute_ctrl1_down_integer_RS2_lane0 = _zz_execute_ctrl1_down_integer_RS2_lane0_1;
  assign when_ExecuteLanePlugin_l196_1 = execute_lane0_bypasser_integer_RS2_sel[0];
  assign execute_lane0_logic_completions_onCtrl_0_port_valid = (((execute_ctrl2_down_LANE_SEL_lane0 && execute_ctrl2_down_isReady) && (! execute_lane0_ctrls_2_downIsCancel)) && execute_ctrl2_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0);
  assign execute_lane0_logic_completions_onCtrl_0_port_payload_uopId = execute_ctrl2_down_Decode_UOP_ID_lane0;
  assign execute_lane0_logic_completions_onCtrl_0_port_payload_trap = execute_ctrl2_down_TRAP_lane0;
  assign execute_lane0_logic_completions_onCtrl_0_port_payload_commit = execute_ctrl2_down_COMMIT_lane0;
  assign execute_lane0_logic_completions_onCtrl_1_port_valid = (((execute_ctrl4_down_LANE_SEL_lane0 && execute_ctrl4_down_isReady) && (! execute_lane0_ctrls_4_downIsCancel)) && execute_ctrl4_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0);
  assign execute_lane0_logic_completions_onCtrl_1_port_payload_uopId = execute_ctrl4_down_Decode_UOP_ID_lane0;
  assign execute_lane0_logic_completions_onCtrl_1_port_payload_trap = execute_ctrl4_down_TRAP_lane0;
  assign execute_lane0_logic_completions_onCtrl_1_port_payload_commit = execute_ctrl4_down_COMMIT_lane0;
  assign execute_lane0_logic_completions_onCtrl_2_port_valid = (((execute_ctrl3_down_LANE_SEL_lane0 && execute_ctrl3_down_isReady) && (! execute_lane0_ctrls_3_downIsCancel)) && execute_ctrl3_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0);
  assign execute_lane0_logic_completions_onCtrl_2_port_payload_uopId = execute_ctrl3_down_Decode_UOP_ID_lane0;
  assign execute_lane0_logic_completions_onCtrl_2_port_payload_trap = execute_ctrl3_down_TRAP_lane0;
  assign execute_lane0_logic_completions_onCtrl_2_port_payload_commit = execute_ctrl3_down_COMMIT_lane0;
  assign execute_lane0_logic_decoding_decodingBits = execute_ctrl1_down_Decode_UOP_lane0;
  assign _zz_execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0 = ((execute_lane0_logic_decoding_decodingBits & 32'h0000004c) == 32'h00000004);
  always @(*) begin
    execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0 = _zz_execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0_1[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_early0_BarrelShifterPlugin_SEL_lane0 = _zz_execute_ctrl1_down_early0_BarrelShifterPlugin_SEL_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_early0_BarrelShifterPlugin_SEL_lane0 = 1'b0;
    end
  end

  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0 = ((execute_lane0_logic_decoding_decodingBits & 32'h00000050) == 32'h00000040);
  always @(*) begin
    execute_ctrl1_down_early0_BranchPlugin_SEL_lane0 = _zz_execute_ctrl1_down_early0_BranchPlugin_SEL_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_early0_BranchPlugin_SEL_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_early0_MulPlugin_SEL_lane0 = _zz_execute_ctrl1_down_early0_MulPlugin_SEL_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_early0_MulPlugin_SEL_lane0 = 1'b0;
    end
  end

  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0 = ((execute_lane0_logic_decoding_decodingBits & 32'h02004064) == 32'h02004020);
  always @(*) begin
    execute_ctrl1_down_early0_DivPlugin_SEL_lane0 = _zz_execute_ctrl1_down_early0_DivPlugin_SEL_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_early0_DivPlugin_SEL_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_early0_EnvPlugin_SEL_lane0 = _zz_execute_ctrl1_down_early0_EnvPlugin_SEL_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_early0_EnvPlugin_SEL_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_MulPlugin_HIGH_lane0 = _zz_execute_ctrl1_down_MulPlugin_HIGH_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_MulPlugin_HIGH_lane0 = 1'b0;
    end
  end

  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0_1 = ((execute_lane0_logic_decoding_decodingBits & 32'h00002050) == 32'h00002050);
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0_2 = ((execute_lane0_logic_decoding_decodingBits & 32'h00001050) == 32'h00001050);
  always @(*) begin
    execute_ctrl1_down_CsrAccessPlugin_SEL_lane0 = _zz_execute_ctrl1_down_CsrAccessPlugin_SEL_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_CsrAccessPlugin_SEL_lane0 = 1'b0;
    end
  end

  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0 = ((execute_lane0_logic_decoding_decodingBits & 32'h00000058) == 32'h0);
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_1 = ((execute_lane0_logic_decoding_decodingBits & 32'h00001050) == 32'h0);
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_2 = ((execute_lane0_logic_decoding_decodingBits & 32'h00002050) == 32'h00002000);
  always @(*) begin
    execute_ctrl1_down_AguPlugin_SEL_lane0 = _zz_execute_ctrl1_down_AguPlugin_SEL_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_AguPlugin_SEL_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_LsuPlugin_logic_FENCE_lane0 = _zz_execute_ctrl1_down_LsuPlugin_logic_FENCE_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_LsuPlugin_logic_FENCE_lane0 = 1'b0;
    end
  end

  assign _zz_execute_ctrl1_down_AguPlugin_LOAD_lane0 = ((execute_lane0_logic_decoding_decodingBits & 32'h00000028) == 32'h0);
  assign _zz_execute_ctrl1_down_BYPASSED_AT_3_lane0 = ((execute_lane0_logic_decoding_decodingBits & 32'h0000000c) == 32'h00000004);
  assign _zz_execute_ctrl1_down_AguPlugin_ATOMIC_lane0 = ((execute_lane0_logic_decoding_decodingBits & 32'h00000028) == 32'h00000028);
  always @(*) begin
    execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0 = _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0 = 1'b0;
    end
  end

  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_1 = ((execute_lane0_logic_decoding_decodingBits & 32'h00007008) == 32'h00001008);
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_2 = ((execute_lane0_logic_decoding_decodingBits & 32'h02000050) == 32'h00000010);
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_3 = ((execute_lane0_logic_decoding_decodingBits & 32'h00003040) == 32'h00000040);
  assign _zz_execute_ctrl1_down_BYPASSED_AT_3_lane0_1 = ((execute_lane0_logic_decoding_decodingBits & 32'h00000030) == 32'h00000010);
  always @(*) begin
    execute_ctrl1_down_COMPLETION_AT_2_lane0 = _zz_execute_ctrl1_down_COMPLETION_AT_2_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_COMPLETION_AT_2_lane0 = 1'b0;
    end
  end

  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_3 = ((execute_lane0_logic_decoding_decodingBits & 32'h02004064) == 32'h02000020);
  always @(*) begin
    execute_ctrl1_down_COMPLETION_AT_4_lane0 = _zz_execute_ctrl1_down_COMPLETION_AT_4_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_COMPLETION_AT_4_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_COMPLETION_AT_3_lane0 = _zz_execute_ctrl1_down_COMPLETION_AT_3_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_COMPLETION_AT_3_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0 = _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_4[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0 = _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_4[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0 = _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0_3[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0 = 1'b0;
    end
  end

  assign _zz_execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0 = ((execute_lane0_logic_decoding_decodingBits & 32'h00006000) == 32'h0);
  assign _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0 = ((execute_lane0_logic_decoding_decodingBits & 32'h00000004) == 32'h00000004);
  assign execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0 = _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0_1[0];
  assign execute_ctrl1_down_early0_IntAluPlugin_ALU_SLTX_lane0 = _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_SLTX_lane0[0];
  assign _zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0 = ((execute_lane0_logic_decoding_decodingBits & 32'h00004000) == 32'h0);
  assign _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0 = ((execute_lane0_logic_decoding_decodingBits & 32'h00001000) == 32'h00001000);
  assign _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1 = {(|{_zz_execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0,{_zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0,_zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0}}),(|{_zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0,{_zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0,((execute_lane0_logic_decoding_decodingBits & 32'h00003000) == 32'h00002000)}})};
  assign _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0 = _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1;
  assign _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2 = _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  assign execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0 = _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2;
  assign _zz_execute_ctrl1_down_BYPASSED_AT_3_lane0_2 = ((execute_lane0_logic_decoding_decodingBits & 32'h00000040) == 32'h00000040);
  assign execute_ctrl1_down_SrcStageables_REVERT_lane0 = _zz_execute_ctrl1_down_SrcStageables_REVERT_lane0[0];
  assign execute_ctrl1_down_SrcStageables_ZERO_lane0 = _zz_execute_ctrl1_down_SrcStageables_ZERO_lane0[0];
  assign execute_ctrl1_down_early0_SrcPlugin_logic_SRC1_CTRL_lane0 = (|_zz_execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0);
  assign execute_ctrl1_down_early0_SrcPlugin_logic_SRC2_CTRL_lane0 = {(|{_zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0,((execute_lane0_logic_decoding_decodingBits & 32'h00000070) == 32'h00000020)}),(|{((execute_lane0_logic_decoding_decodingBits & 32'h00000050) == 32'h0),((execute_lane0_logic_decoding_decodingBits & 32'h00000024) == 32'h0)})};
  assign _zz_execute_ctrl1_down_RsUnsignedPlugin_IS_W_lane0 = ((execute_lane0_logic_decoding_decodingBits & 32'h00000008) == 32'h00000008);
  assign execute_ctrl1_down_lane0_IntFormatPlugin_logic_SIGNED_lane0 = _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_SIGNED_lane0[0];
  assign _zz_execute_ctrl1_down_AguPlugin_STORE_lane0 = ((execute_lane0_logic_decoding_decodingBits & 32'h10000020) == 32'h00000020);
  assign execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0 = {(|{((execute_lane0_logic_decoding_decodingBits & _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0) == 32'h00000010),{(_zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0_1 == _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0_2),{_zz_execute_ctrl1_down_AguPlugin_STORE_lane0,_zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0_3}}}),(|{((execute_lane0_logic_decoding_decodingBits & _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0_4) == 32'h00000010),{(_zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0_5 == _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0_6),{_zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0_7,_zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0_8}}})};
  assign execute_ctrl1_down_BYPASSED_AT_2_lane0 = _zz_execute_ctrl1_down_BYPASSED_AT_2_lane0[0];
  assign execute_ctrl1_down_BYPASSED_AT_3_lane0 = _zz_execute_ctrl1_down_BYPASSED_AT_3_lane0_3[0];
  assign execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane0 = _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane0[0];
  assign execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane0 = _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane0[0];
  assign execute_ctrl1_down_SrcStageables_UNSIGNED_lane0 = _zz_execute_ctrl1_down_SrcStageables_UNSIGNED_lane0[0];
  assign execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0 = _zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0_1[0];
  assign execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane0 = _zz_execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane0[0];
  assign execute_ctrl1_down_BarrelShifterPlugin_IS_W_lane0 = _zz_execute_ctrl1_down_BarrelShifterPlugin_IS_W_lane0[0];
  assign execute_ctrl1_down_BarrelShifterPlugin_IS_W_RIGHT_lane0 = _zz_execute_ctrl1_down_BarrelShifterPlugin_IS_W_RIGHT_lane0[0];
  assign _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_1 = {(|_zz_execute_ctrl1_down_BYPASSED_AT_3_lane0),(|_zz_execute_ctrl1_down_RsUnsignedPlugin_IS_W_lane0)};
  assign _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0 = _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_1;
  assign _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_2 = _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0;
  assign execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0 = _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_2;
  assign execute_ctrl1_down_RsUnsignedPlugin_RS1_SIGNED_lane0 = _zz_execute_ctrl1_down_RsUnsignedPlugin_RS1_SIGNED_lane0[0];
  assign execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0 = _zz_execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0_1[0];
  assign _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0 = ((execute_lane0_logic_decoding_decodingBits & 32'h00002000) == 32'h00002000);
  assign execute_ctrl1_down_DivPlugin_REM_lane0 = _zz_execute_ctrl1_down_DivPlugin_REM_lane0[0];
  assign execute_ctrl1_down_RsUnsignedPlugin_IS_W_lane0 = _zz_execute_ctrl1_down_RsUnsignedPlugin_IS_W_lane0_1[0];
  assign execute_ctrl1_down_CsrAccessPlugin_CSR_IMM_lane0 = _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_IMM_lane0[0];
  assign execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0 = _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0_1[0];
  assign execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0 = _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0_1[0];
  assign execute_ctrl1_down_AguPlugin_LOAD_lane0 = _zz_execute_ctrl1_down_AguPlugin_LOAD_lane0_1[0];
  assign execute_ctrl1_down_AguPlugin_STORE_lane0 = _zz_execute_ctrl1_down_AguPlugin_STORE_lane0_1[0];
  assign execute_ctrl1_down_AguPlugin_ATOMIC_lane0 = _zz_execute_ctrl1_down_AguPlugin_ATOMIC_lane0_1[0];
  assign execute_ctrl1_down_AguPlugin_FLOAT_lane0 = _zz_execute_ctrl1_down_AguPlugin_FLOAT_lane0[0];
  assign execute_ctrl1_down_AguPlugin_CLEAN_lane0 = _zz_execute_ctrl1_down_AguPlugin_CLEAN_lane0[0];
  assign execute_ctrl1_down_AguPlugin_INVALIDATE_lane0 = _zz_execute_ctrl1_down_AguPlugin_INVALIDATE_lane0[0];
  assign execute_ctrl1_down_LsuPlugin_logic_LSU_PREFETCH_lane0 = _zz_execute_ctrl1_down_LsuPlugin_logic_LSU_PREFETCH_lane0[0];
  assign _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0 = ((execute_lane0_logic_decoding_decodingBits & 32'h00000040) == 32'h0);
  assign _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2 = {(|{((execute_lane0_logic_decoding_decodingBits & _zz__zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2) == 32'h02000000),((execute_lane0_logic_decoding_decodingBits & _zz__zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_1) == 32'h10000000)}),{(|{_zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0,(_zz__zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_2 == _zz__zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_3)}),(|{_zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0,{_zz__zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_4,_zz__zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_5}})}};
  assign _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1 = _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2;
  assign _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_3 = _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1;
  assign execute_ctrl1_down_early0_EnvPlugin_OP_lane0 = _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_3;
  assign when_ExecuteLanePlugin_l306 = (|{(early0_EnvPlugin_logic_flushPort_valid && 1'b1),{(CsrAccessPlugin_logic_flushPort_valid && 1'b1),{(early0_BranchPlugin_logic_flushPort_valid && 1'b1),(LsuPlugin_logic_flushPort_valid && 1'b1)}}});
  assign execute_lane0_ctrls_0_downIsCancel = 1'b0;
  assign execute_lane0_ctrls_0_upIsCancel = when_ExecuteLanePlugin_l306;
  assign when_ExecuteLanePlugin_l306_1 = (|{(early0_EnvPlugin_logic_flushPort_valid && 1'b1),{(CsrAccessPlugin_logic_flushPort_valid && 1'b1),{(early0_BranchPlugin_logic_flushPort_valid && 1'b1),(LsuPlugin_logic_flushPort_valid && 1'b1)}}});
  assign execute_lane0_ctrls_1_downIsCancel = 1'b0;
  assign execute_lane0_ctrls_1_upIsCancel = when_ExecuteLanePlugin_l306_1;
  assign when_ExecuteLanePlugin_l306_2 = (|{((early0_EnvPlugin_logic_flushPort_valid && 1'b1) && (1'b0 || (1'b1 && early0_EnvPlugin_logic_flushPort_payload_self))),{((CsrAccessPlugin_logic_flushPort_valid && 1'b1) && (1'b0 || (_zz_when_ExecuteLanePlugin_l306_2 && CsrAccessPlugin_logic_flushPort_payload_self))),{((early0_BranchPlugin_logic_flushPort_valid && _zz_when_ExecuteLanePlugin_l306_2_1) && (_zz_when_ExecuteLanePlugin_l306_2_2 || _zz_when_ExecuteLanePlugin_l306_2_3)),(LsuPlugin_logic_flushPort_valid && 1'b1)}}});
  assign execute_lane0_ctrls_2_downIsCancel = 1'b0;
  assign execute_lane0_ctrls_2_upIsCancel = when_ExecuteLanePlugin_l306_2;
  assign when_ExecuteLanePlugin_l306_3 = (|(LsuPlugin_logic_flushPort_valid && 1'b1));
  assign execute_lane0_ctrls_3_downIsCancel = 1'b0;
  assign execute_lane0_ctrls_3_upIsCancel = when_ExecuteLanePlugin_l306_3;
  assign when_ExecuteLanePlugin_l306_4 = (|((LsuPlugin_logic_flushPort_valid && 1'b1) && (1'b0 || (1'b1 && LsuPlugin_logic_flushPort_payload_self))));
  assign execute_lane0_ctrls_4_downIsCancel = 1'b0;
  assign execute_lane0_ctrls_4_upIsCancel = when_ExecuteLanePlugin_l306_4;
  assign execute_lane0_ctrls_5_downIsCancel = 1'b0;
  assign execute_lane0_ctrls_5_upIsCancel = 1'b0;
  assign execute_lane0_logic_trapPending[0] = (|{((execute_ctrl4_up_LANE_SEL_lane0 && 1'b1) && execute_ctrl4_down_TRAP_lane0),{((execute_ctrl3_up_LANE_SEL_lane0 && 1'b1) && execute_ctrl3_down_TRAP_lane0),{((execute_ctrl2_up_LANE_SEL_lane0 && 1'b1) && execute_ctrl2_down_TRAP_lane0),((execute_ctrl1_up_LANE_SEL_lane0 && 1'b1) && execute_ctrl1_down_TRAP_lane0)}}});
  assign execute_ctrl2_up_COMMIT_lane0 = (! execute_ctrl2_up_TRAP_lane0);
  assign WhiteboxerPlugin_logic_csr_access_valid = CsrAccessPlugin_logic_fsm_interface_fire;
  assign WhiteboxerPlugin_logic_csr_access_payload_uopId = CsrAccessPlugin_logic_fsm_interface_uopId;
  assign WhiteboxerPlugin_logic_csr_access_payload_address = _zz_WhiteboxerPlugin_logic_csr_access_payload_address[31 : 20];
  assign WhiteboxerPlugin_logic_csr_access_payload_write = CsrAccessPlugin_logic_fsm_interface_onWriteBits;
  assign WhiteboxerPlugin_logic_csr_access_payload_read = CsrAccessPlugin_logic_fsm_interface_csrValue;
  assign WhiteboxerPlugin_logic_csr_access_payload_writeDone = CsrAccessPlugin_logic_fsm_interface_write;
  assign WhiteboxerPlugin_logic_csr_access_payload_readDone = CsrAccessPlugin_logic_fsm_interface_read;
  assign WhiteboxerPlugin_logic_csr_port_valid = WhiteboxerPlugin_logic_csr_access_valid;
  assign WhiteboxerPlugin_logic_csr_port_payload_uopId = WhiteboxerPlugin_logic_csr_access_payload_uopId;
  assign WhiteboxerPlugin_logic_csr_port_payload_address = WhiteboxerPlugin_logic_csr_access_payload_address;
  assign WhiteboxerPlugin_logic_csr_port_payload_write = WhiteboxerPlugin_logic_csr_access_payload_write;
  assign WhiteboxerPlugin_logic_csr_port_payload_read = WhiteboxerPlugin_logic_csr_access_payload_read;
  assign WhiteboxerPlugin_logic_csr_port_payload_writeDone = WhiteboxerPlugin_logic_csr_access_payload_writeDone;
  assign WhiteboxerPlugin_logic_csr_port_payload_readDone = WhiteboxerPlugin_logic_csr_access_payload_readDone;
  assign WhiteboxerPlugin_logic_rfWrites_ports_0_valid = lane0_integer_WriteBackPlugin_logic_stages_0_write_valid;
  assign WhiteboxerPlugin_logic_rfWrites_ports_0_payload_uopId = lane0_integer_WriteBackPlugin_logic_stages_0_write_payload_uopId;
  assign WhiteboxerPlugin_logic_rfWrites_ports_0_payload_data = lane0_integer_WriteBackPlugin_logic_stages_0_write_payload_data;
  assign WhiteboxerPlugin_logic_rfWrites_ports_1_valid = lane0_integer_WriteBackPlugin_logic_stages_1_write_valid;
  assign WhiteboxerPlugin_logic_rfWrites_ports_1_payload_uopId = lane0_integer_WriteBackPlugin_logic_stages_1_write_payload_uopId;
  assign WhiteboxerPlugin_logic_rfWrites_ports_1_payload_data = lane0_integer_WriteBackPlugin_logic_stages_1_write_payload_data;
  assign WhiteboxerPlugin_logic_rfWrites_ports_2_valid = lane0_integer_WriteBackPlugin_logic_stages_2_write_valid;
  assign WhiteboxerPlugin_logic_rfWrites_ports_2_payload_uopId = lane0_integer_WriteBackPlugin_logic_stages_2_write_payload_uopId;
  assign WhiteboxerPlugin_logic_rfWrites_ports_2_payload_data = lane0_integer_WriteBackPlugin_logic_stages_2_write_payload_data;
  assign WhiteboxerPlugin_logic_completions_ports_0_valid = DecoderPlugin_logic_laneLogic_0_completionPort_valid;
  assign WhiteboxerPlugin_logic_completions_ports_0_payload_uopId = DecoderPlugin_logic_laneLogic_0_completionPort_payload_uopId;
  assign WhiteboxerPlugin_logic_completions_ports_0_payload_trap = DecoderPlugin_logic_laneLogic_0_completionPort_payload_trap;
  assign WhiteboxerPlugin_logic_completions_ports_0_payload_commit = DecoderPlugin_logic_laneLogic_0_completionPort_payload_commit;
  assign WhiteboxerPlugin_logic_completions_ports_1_valid = execute_lane0_logic_completions_onCtrl_0_port_valid;
  assign WhiteboxerPlugin_logic_completions_ports_1_payload_uopId = execute_lane0_logic_completions_onCtrl_0_port_payload_uopId;
  assign WhiteboxerPlugin_logic_completions_ports_1_payload_trap = execute_lane0_logic_completions_onCtrl_0_port_payload_trap;
  assign WhiteboxerPlugin_logic_completions_ports_1_payload_commit = execute_lane0_logic_completions_onCtrl_0_port_payload_commit;
  assign WhiteboxerPlugin_logic_completions_ports_2_valid = execute_lane0_logic_completions_onCtrl_1_port_valid;
  assign WhiteboxerPlugin_logic_completions_ports_2_payload_uopId = execute_lane0_logic_completions_onCtrl_1_port_payload_uopId;
  assign WhiteboxerPlugin_logic_completions_ports_2_payload_trap = execute_lane0_logic_completions_onCtrl_1_port_payload_trap;
  assign WhiteboxerPlugin_logic_completions_ports_2_payload_commit = execute_lane0_logic_completions_onCtrl_1_port_payload_commit;
  assign WhiteboxerPlugin_logic_completions_ports_3_valid = execute_lane0_logic_completions_onCtrl_2_port_valid;
  assign WhiteboxerPlugin_logic_completions_ports_3_payload_uopId = execute_lane0_logic_completions_onCtrl_2_port_payload_uopId;
  assign WhiteboxerPlugin_logic_completions_ports_3_payload_trap = execute_lane0_logic_completions_onCtrl_2_port_payload_trap;
  assign WhiteboxerPlugin_logic_completions_ports_3_payload_commit = execute_lane0_logic_completions_onCtrl_2_port_payload_commit;
  assign WhiteboxerPlugin_logic_commits_ports_0_oh_0 = ((((execute_ctrl4_down_LANE_SEL_lane0 && execute_ctrl4_down_isReady) && (! execute_lane0_ctrls_4_downIsCancel)) && execute_ctrl4_down_COMMIT_lane0) && 1'b1);
  assign WhiteboxerPlugin_logic_commits_ports_0_valid = (|WhiteboxerPlugin_logic_commits_ports_0_oh_0);
  assign WhiteboxerPlugin_logic_commits_ports_0_pc = (WhiteboxerPlugin_logic_commits_ports_0_oh_0 ? execute_ctrl4_down_PC_lane0 : 39'h0);
  assign WhiteboxerPlugin_logic_commits_ports_0_uop = (WhiteboxerPlugin_logic_commits_ports_0_oh_0 ? execute_ctrl4_down_Decode_UOP_lane0 : 32'h0);
  assign WhiteboxerPlugin_logic_reschedules_flushes_0_valid = BtbPlugin_logic_flushPort_valid;
  assign WhiteboxerPlugin_logic_reschedules_flushes_0_payload_self = BtbPlugin_logic_flushPort_payload_self;
  assign WhiteboxerPlugin_logic_reschedules_flushes_1_valid = LsuPlugin_logic_flushPort_valid;
  assign WhiteboxerPlugin_logic_reschedules_flushes_1_payload_uopId = LsuPlugin_logic_flushPort_payload_uopId;
  assign WhiteboxerPlugin_logic_reschedules_flushes_1_payload_self = LsuPlugin_logic_flushPort_payload_self;
  assign WhiteboxerPlugin_logic_reschedules_flushes_2_valid = early0_BranchPlugin_logic_flushPort_valid;
  assign WhiteboxerPlugin_logic_reschedules_flushes_2_payload_uopId = early0_BranchPlugin_logic_flushPort_payload_uopId;
  assign WhiteboxerPlugin_logic_reschedules_flushes_2_payload_self = early0_BranchPlugin_logic_flushPort_payload_self;
  assign WhiteboxerPlugin_logic_reschedules_flushes_3_valid = CsrAccessPlugin_logic_flushPort_valid;
  assign WhiteboxerPlugin_logic_reschedules_flushes_3_payload_uopId = CsrAccessPlugin_logic_flushPort_payload_uopId;
  assign WhiteboxerPlugin_logic_reschedules_flushes_3_payload_self = CsrAccessPlugin_logic_flushPort_payload_self;
  assign WhiteboxerPlugin_logic_reschedules_flushes_4_valid = early0_EnvPlugin_logic_flushPort_valid;
  assign WhiteboxerPlugin_logic_reschedules_flushes_4_payload_uopId = early0_EnvPlugin_logic_flushPort_payload_uopId;
  assign WhiteboxerPlugin_logic_reschedules_flushes_4_payload_self = early0_EnvPlugin_logic_flushPort_payload_self;
  assign WhiteboxerPlugin_logic_reschedules_flushes_5_valid = DecoderPlugin_logic_laneLogic_0_flushPort_valid;
  assign WhiteboxerPlugin_logic_reschedules_flushes_5_payload_uopId = DecoderPlugin_logic_laneLogic_0_flushPort_payload_uopId;
  assign WhiteboxerPlugin_logic_reschedules_flushes_5_payload_self = DecoderPlugin_logic_laneLogic_0_flushPort_payload_self;
  assign early0_BranchPlugin_logic_jumpLogic_learn_asFlow_valid = early0_BranchPlugin_logic_jumpLogic_learn_valid;
  assign early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_pcOnLastSlice = early0_BranchPlugin_logic_jumpLogic_learn_payload_pcOnLastSlice;
  assign early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_pcTarget = early0_BranchPlugin_logic_jumpLogic_learn_payload_pcTarget;
  assign early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_taken = early0_BranchPlugin_logic_jumpLogic_learn_payload_taken;
  assign early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_isBranch = early0_BranchPlugin_logic_jumpLogic_learn_payload_isBranch;
  assign early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_isPush = early0_BranchPlugin_logic_jumpLogic_learn_payload_isPush;
  assign early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_isPop = early0_BranchPlugin_logic_jumpLogic_learn_payload_isPop;
  assign early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_wasWrong = early0_BranchPlugin_logic_jumpLogic_learn_payload_wasWrong;
  assign early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_badPredictedTarget = early0_BranchPlugin_logic_jumpLogic_learn_payload_badPredictedTarget;
  assign early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_history = early0_BranchPlugin_logic_jumpLogic_learn_payload_history;
  assign early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_uopId = early0_BranchPlugin_logic_jumpLogic_learn_payload_uopId;
  assign early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 = early0_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  assign early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_1 = early0_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  assign WhiteboxerPlugin_logic_prediction_learns_0_valid = early0_BranchPlugin_logic_jumpLogic_learn_asFlow_valid;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_pcOnLastSlice = early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_pcOnLastSlice;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_pcTarget = early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_pcTarget;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_taken = early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_taken;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_isBranch = early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_isBranch;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_isPush = early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_isPush;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_isPop = early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_isPop;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_wasWrong = early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_wasWrong;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_badPredictedTarget = early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_badPredictedTarget;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_history = early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_history;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_uopId = early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_uopId;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 = early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_1 = early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  assign WhiteboxerPlugin_logic_loadExecute_fire = (((((((execute_ctrl4_down_LANE_SEL_lane0 && execute_ctrl4_down_isReady) && (! execute_lane0_ctrls_4_downIsCancel)) && execute_ctrl4_down_AguPlugin_SEL_lane0) && execute_ctrl4_down_AguPlugin_LOAD_lane0) && (! execute_ctrl4_down_LsuPlugin_logic_LSU_PREFETCH_lane0)) && (! execute_ctrl4_down_TRAP_lane0)) && (! execute_ctrl4_down_LsuPlugin_logic_onPma_IO_lane0));
  assign WhiteboxerPlugin_logic_loadExecute_uopId = execute_ctrl4_down_Decode_UOP_ID_lane0;
  assign WhiteboxerPlugin_logic_loadExecute_size = execute_ctrl4_down_AguPlugin_SIZE_lane0;
  assign WhiteboxerPlugin_logic_loadExecute_address = execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0;
  assign WhiteboxerPlugin_logic_loadExecute_data = lane0_IntFormatPlugin_logic_stages_1_wb_payload;
  assign WhiteboxerPlugin_logic_storeCommit_fire = LsuPlugin_logic_onWb_storeFire;
  assign WhiteboxerPlugin_logic_storeCommit_uopId = execute_ctrl4_down_Decode_UOP_ID_lane0;
  assign WhiteboxerPlugin_logic_storeCommit_size = execute_ctrl4_down_AguPlugin_SIZE_lane0;
  assign WhiteboxerPlugin_logic_storeCommit_address = execute_ctrl4_down_MMU_TRANSLATED_lane0;
  assign WhiteboxerPlugin_logic_storeCommit_data = execute_ctrl4_down_LsuL1_WRITE_DATA_lane0;
  assign WhiteboxerPlugin_logic_storeCommit_storeId = execute_ctrl4_down_Decode_STORE_ID_lane0;
  assign WhiteboxerPlugin_logic_storeCommit_amo = 1'b0;
  assign WhiteboxerPlugin_logic_storeConditional_fire = (((((execute_ctrl4_down_LANE_SEL_lane0 && execute_ctrl4_down_isReady) && (! execute_lane0_ctrls_4_downIsCancel)) && execute_ctrl4_down_AguPlugin_SEL_lane0) && (execute_ctrl4_down_AguPlugin_ATOMIC_lane0 && (! execute_ctrl4_down_AguPlugin_LOAD_lane0))) && (! execute_ctrl4_down_TRAP_lane0));
  assign WhiteboxerPlugin_logic_storeConditional_uopId = execute_ctrl4_down_Decode_UOP_ID_lane0;
  assign WhiteboxerPlugin_logic_storeConditional_miss = execute_ctrl4_down_LsuPlugin_logic_onCtrl_SC_MISS_lane0;
  assign WhiteboxerPlugin_logic_storeBroadcast_fire = LsuPlugin_logic_onWb_storeBroadcast;
  assign WhiteboxerPlugin_logic_storeBroadcast_storeId = execute_ctrl4_down_Decode_STORE_ID_lane0;
  assign integer_RegFilePlugin_logic_writeMerges_0_bus_valid = (|lane0_integer_WriteBackPlugin_logic_write_port_valid);
  assign integer_RegFilePlugin_logic_writeMerges_0_bus_address = lane0_integer_WriteBackPlugin_logic_write_port_address;
  assign integer_RegFilePlugin_logic_writeMerges_0_bus_data = lane0_integer_WriteBackPlugin_logic_write_port_data;
  assign integer_RegFilePlugin_logic_writeMerges_0_bus_uopId = lane0_integer_WriteBackPlugin_logic_write_port_uopId;
  assign execute_lane0_bypasser_integer_RS1_port_data = integer_RegFilePlugin_logic_regfile_fpga_io_reads_0_data;
  assign execute_lane0_bypasser_integer_RS2_port_data = integer_RegFilePlugin_logic_regfile_fpga_io_reads_1_data;
  always @(*) begin
    integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_valid = integer_RegFilePlugin_logic_writeMerges_0_bus_valid;
    if(when_RegFilePlugin_l132) begin
      integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_valid = 1'b1;
    end
  end

  always @(*) begin
    integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_address = integer_RegFilePlugin_logic_writeMerges_0_bus_address;
    if(when_RegFilePlugin_l132) begin
      integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_address = integer_RegFilePlugin_logic_initalizer_counter[4:0];
    end
  end

  always @(*) begin
    integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_data = integer_RegFilePlugin_logic_writeMerges_0_bus_data;
    if(when_RegFilePlugin_l132) begin
      integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_data = 64'h0;
    end
  end

  assign integer_RegFilePlugin_logic_initalizer_done = integer_RegFilePlugin_logic_initalizer_counter[5];
  assign when_RegFilePlugin_l132 = (! integer_RegFilePlugin_logic_initalizer_done);
  assign integer_write_0_valid = integer_RegFilePlugin_logic_writeMerges_0_bus_valid;
  assign integer_write_0_address = integer_RegFilePlugin_logic_writeMerges_0_bus_address;
  assign integer_write_0_data = integer_RegFilePlugin_logic_writeMerges_0_bus_data;
  assign integer_write_0_uopId = integer_RegFilePlugin_logic_writeMerges_0_bus_uopId;
  assign execute_freeze_valid = (|{CsrAccessPlugin_logic_fsm_inject_freeze,{LsuPlugin_logic_onCtrl_rva_freezeIt,{LsuPlugin_logic_onCtrl_io_freezeIt,{early0_DivPlugin_logic_processing_freeze,((execute_ctrl4_up_LANE_SEL_lane0 && execute_ctrl4_down_MulPlugin_HIGH_lane0) && (! early0_MulPlugin_logic_writeback_buffer_valid))}}}});
  assign execute_ctrl5_down_ready = (! execute_freeze_valid);
  assign TrapPlugin_logic_initHold = (|{(! CsrRamPlugin_logic_flush_done),{((! LsuL1Plugin_logic_initializer_done) || 1'b0),{(! integer_RegFilePlugin_logic_initalizer_done),{(FetchL1Plugin_logic_invalidate_firstEver || 1'b0),{1'b0,1'b0}}}}});
  assign WhiteboxerPlugin_logic_wfi = TrapPlugin_logic_harts_0_trap_fsm_wfi;
  assign WhiteboxerPlugin_logic_perf_executeFreezed = execute_freeze_valid;
  assign WhiteboxerPlugin_logic_perf_dispatchHazards = (|(DispatchPlugin_logic_candidates_0_ctx_valid && (! DispatchPlugin_logic_candidates_0_fire)));
  assign WhiteboxerPlugin_logic_perf_candidatesCount = _zz_WhiteboxerPlugin_logic_perf_candidatesCount;
  assign WhiteboxerPlugin_logic_perf_dispatchFeedCount = _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCount;
  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter = 1'b0;
    if(WhiteboxerPlugin_logic_perf_executeFreezed) begin
      _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter = 1'b1;
    end
  end

  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_1 = (_zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_2 + _zz__zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_1);
    if(1'b0) begin
      _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_1 = 60'h0;
    end
  end

  assign WhiteboxerPlugin_logic_perf_executeFreezedCounter = _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_2;
  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter = 1'b0;
    if(WhiteboxerPlugin_logic_perf_dispatchHazards) begin
      _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter = 1'b1;
    end
  end

  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_1 = (_zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_2 + _zz__zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_1);
    if(1'b0) begin
      _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_1 = 60'h0;
    end
  end

  assign WhiteboxerPlugin_logic_perf_dispatchHazardsCounter = _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_2;
  assign when_Utils_l598 = (WhiteboxerPlugin_logic_perf_candidatesCount == 1'b0);
  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0 = 1'b0;
    if(when_Utils_l598) begin
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0 = 1'b1;
    end
  end

  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_1 = (_zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_2 + _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_1);
    if(1'b0) begin
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_1 = 60'h0;
    end
  end

  assign WhiteboxerPlugin_logic_perf_candidatesCountCounters_0 = _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_2;
  assign when_Utils_l598_1 = (WhiteboxerPlugin_logic_perf_candidatesCount == 1'b1);
  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1 = 1'b0;
    if(when_Utils_l598_1) begin
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1 = 1'b1;
    end
  end

  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_1 = (_zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_2 + _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_1);
    if(1'b0) begin
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_1 = 60'h0;
    end
  end

  assign WhiteboxerPlugin_logic_perf_candidatesCountCounters_1 = _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_2;
  assign when_Utils_l598_2 = (WhiteboxerPlugin_logic_perf_dispatchFeedCount == 1'b0);
  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0 = 1'b0;
    if(when_Utils_l598_2) begin
      _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0 = 1'b1;
    end
  end

  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_1 = (_zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_2 + _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_1);
    if(1'b0) begin
      _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_1 = 60'h0;
    end
  end

  assign WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0 = _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_2;
  assign when_Utils_l598_3 = (WhiteboxerPlugin_logic_perf_dispatchFeedCount == 1'b1);
  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1 = 1'b0;
    if(when_Utils_l598_3) begin
      _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1 = 1'b1;
    end
  end

  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_1 = (_zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_2 + _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_1);
    if(1'b0) begin
      _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_1 = 60'h0;
    end
  end

  assign WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1 = _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_2;
  assign WhiteboxerPlugin_logic_trap_ports_0_valid = TrapPlugin_logic_harts_0_trap_whitebox_trap;
  assign WhiteboxerPlugin_logic_trap_ports_0_interrupt = TrapPlugin_logic_harts_0_trap_whitebox_interrupt;
  assign WhiteboxerPlugin_logic_trap_ports_0_cause = TrapPlugin_logic_harts_0_trap_whitebox_code;
  assign fetch_logic_ctrls_2_up_forgetOne = (|fetch_logic_ctrls_2_forgetsSingleRequest_FetchPipelinePlugin_l50);
  assign fetch_logic_ctrls_2_up_cancel = (|fetch_logic_flushes_1_doIt);
  assign fetch_logic_ctrls_1_up_forgetOne = (|fetch_logic_ctrls_1_throwWhen_FetchPipelinePlugin_l48);
  assign fetch_logic_ctrls_1_up_cancel = (|fetch_logic_ctrls_1_throwWhen_FetchPipelinePlugin_l48);
  assign fetch_logic_ctrls_0_down_ready = fetch_logic_ctrls_1_up_ready;
  assign fetch_logic_ctrls_1_down_ready = fetch_logic_ctrls_2_up_ready;
  always @(*) begin
    fetch_logic_ctrls_0_down_valid = fetch_logic_ctrls_0_up_valid;
    if(when_CtrlLink_l191) begin
      fetch_logic_ctrls_0_down_valid = 1'b0;
    end
  end

  always @(*) begin
    fetch_logic_ctrls_0_up_ready = fetch_logic_ctrls_0_down_isReady;
    if(when_CtrlLink_l191) begin
      fetch_logic_ctrls_0_up_ready = 1'b0;
    end
  end

  assign when_CtrlLink_l191 = (|{fetch_logic_ctrls_0_haltRequest_PcPlugin_l133,{fetch_logic_ctrls_0_haltRequest_BtbPlugin_l200,{fetch_logic_ctrls_0_haltRequest_FetchL1Plugin_l297,fetch_logic_ctrls_0_haltRequest_FetchL1Plugin_l217}}});
  assign fetch_logic_ctrls_0_down_Fetch_WORD_PC = fetch_logic_ctrls_0_up_Fetch_WORD_PC;
  assign fetch_logic_ctrls_0_down_Fetch_PC_FAULT = fetch_logic_ctrls_0_up_Fetch_PC_FAULT;
  assign fetch_logic_ctrls_0_down_Fetch_ID = fetch_logic_ctrls_0_up_Fetch_ID;
  always @(*) begin
    fetch_logic_ctrls_1_down_valid = fetch_logic_ctrls_1_up_valid;
    if(when_CtrlLink_l198) begin
      fetch_logic_ctrls_1_down_valid = 1'b0;
    end
  end

  assign fetch_logic_ctrls_1_up_ready = fetch_logic_ctrls_1_down_isReady;
  assign when_CtrlLink_l198 = (|fetch_logic_ctrls_1_throwWhen_FetchPipelinePlugin_l48);
  assign fetch_logic_ctrls_1_down_Fetch_WORD_PC = fetch_logic_ctrls_1_up_Fetch_WORD_PC;
  assign fetch_logic_ctrls_1_down_Fetch_PC_FAULT = fetch_logic_ctrls_1_up_Fetch_PC_FAULT;
  assign fetch_logic_ctrls_1_down_Fetch_ID = fetch_logic_ctrls_1_up_Fetch_ID;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_VALID = fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_PLRU_BYPASS_VALID;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_0 = fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_0;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE = fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_TAGS_UPDATE;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE_ADDRESS = fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_TAGS_UPDATE_ADDRESS;
  assign fetch_logic_ctrls_1_down_GSharePlugin_logic_HASH = fetch_logic_ctrls_1_up_GSharePlugin_logic_HASH;
  assign fetch_logic_ctrls_1_down_Prediction_BRANCH_HISTORY = fetch_logic_ctrls_1_up_Prediction_BRANCH_HISTORY;
  assign fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_valid = fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_valid;
  assign fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_address = fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_address;
  assign fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_data_0 = fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_data_0;
  assign fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_data_1 = fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_data_1;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_PERM_OK = fetch_logic_ctrls_1_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_PERM_OK;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_PERM_OK = fetch_logic_ctrls_1_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_PERM_OK;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_PERM_OK = fetch_logic_ctrls_1_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_PERM_OK;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_PERM_OK = fetch_logic_ctrls_1_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_PERM_OK;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_NEED_HIT = fetch_logic_ctrls_1_up_FetchL1Plugin_logic_pmpPort_logic_NEED_HIT;
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_readCmd_HAZARDS = fetch_logic_ctrls_1_up_BtbPlugin_logic_readCmd_HAZARDS;
  assign fetch_logic_ctrls_2_down_valid = fetch_logic_ctrls_2_up_valid;
  assign fetch_logic_ctrls_2_up_ready = fetch_logic_ctrls_2_down_isReady;
  assign fetch_logic_ctrls_2_down_Fetch_WORD_PC = fetch_logic_ctrls_2_up_Fetch_WORD_PC;
  assign fetch_logic_ctrls_2_down_Fetch_PC_FAULT = fetch_logic_ctrls_2_up_Fetch_PC_FAULT;
  assign fetch_logic_ctrls_2_down_Fetch_ID = fetch_logic_ctrls_2_up_Fetch_ID;
  assign fetch_logic_ctrls_2_down_Prediction_BRANCH_HISTORY = fetch_logic_ctrls_2_up_Prediction_BRANCH_HISTORY;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_PERM_OK = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_PERM_OK;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_PERM_OK = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_PERM_OK;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_PERM_OK = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_PERM_OK;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_PERM_OK = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_PERM_OK;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_NEED_HIT = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_pmpPort_logic_NEED_HIT;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_0_loaded = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_0_loaded;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_0_error = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_0_error;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_0_address = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_0_address;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_1_loaded = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_1_loaded;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_1_error = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_1_error;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_1_address = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_1_address;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_PLRU_BYPASSED_0 = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_PLRU_BYPASSED_0;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_BANKS_MUXES_0 = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_BANKS_MUXES_0;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_BANKS_MUXES_1 = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_BANKS_MUXES_1;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_HAZARD = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_HAZARD;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_0 = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_HITS_0;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_1 = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_HITS_1;
  assign fetch_logic_ctrls_2_down_MMU_BYPASS_TRANSLATION = fetch_logic_ctrls_2_up_MMU_BYPASS_TRANSLATION;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HIT = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_HIT;
  assign fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_0 = fetch_logic_ctrls_2_up_GSharePlugin_GSHARE_COUNTER_0;
  assign fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_1 = fetch_logic_ctrls_2_up_GSharePlugin_GSHARE_COUNTER_1;
  assign fetch_logic_ctrls_2_down_MMU_TRANSLATED = fetch_logic_ctrls_2_up_MMU_TRANSLATED;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_napot_HIT = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_napot_HIT;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_tor_BIGGER = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_tor_BIGGER;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_napot_HIT = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_napot_HIT;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_tor_BIGGER = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_tor_BIGGER;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_napot_HIT = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_napot_HIT;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_tor_BIGGER = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_tor_BIGGER;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_napot_HIT = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_napot_HIT;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_tor_BIGGER = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_tor_BIGGER;
  assign fetch_logic_ctrls_2_down_Prediction_WORD_JUMPED = fetch_logic_ctrls_2_up_Prediction_WORD_JUMPED;
  assign fetch_logic_ctrls_2_down_Prediction_WORD_JUMP_SLICE = fetch_logic_ctrls_2_up_Prediction_WORD_JUMP_SLICE;
  assign fetch_logic_ctrls_2_down_Prediction_WORD_JUMP_PC = fetch_logic_ctrls_2_up_Prediction_WORD_JUMP_PC;
  assign fetch_logic_ctrls_2_down_Prediction_WORD_SLICES_BRANCH = fetch_logic_ctrls_2_up_Prediction_WORD_SLICES_BRANCH;
  assign fetch_logic_ctrls_2_down_Prediction_WORD_SLICES_TAKEN = fetch_logic_ctrls_2_up_Prediction_WORD_SLICES_TAKEN;
  assign fetch_logic_ctrls_2_down_MMU_HAZARD = fetch_logic_ctrls_2_up_MMU_HAZARD;
  assign fetch_logic_ctrls_2_down_MMU_REFILL = fetch_logic_ctrls_2_up_MMU_REFILL;
  assign fetch_logic_ctrls_2_down_MMU_ALLOW_EXECUTE = fetch_logic_ctrls_2_up_MMU_ALLOW_EXECUTE;
  assign fetch_logic_ctrls_2_down_MMU_PAGE_FAULT = fetch_logic_ctrls_2_up_MMU_PAGE_FAULT;
  assign fetch_logic_ctrls_2_down_MMU_ACCESS_FAULT = fetch_logic_ctrls_2_up_MMU_ACCESS_FAULT;
  always @(*) begin
    decode_ctrls_0_down_ready = decode_ctrls_1_up_ready;
    if(when_StageLink_l71) begin
      decode_ctrls_0_down_ready = 1'b1;
    end
  end

  assign when_StageLink_l71 = (! decode_ctrls_1_up_isValid);
  assign when_DecodePipelinePlugin_l70 = ((! decode_ctrls_1_up_isReady) && decode_ctrls_1_lane0_upIsCancel);
  assign decode_ctrls_0_down_valid = decode_ctrls_0_up_valid;
  assign decode_ctrls_0_up_ready = decode_ctrls_0_down_isReady;
  assign decode_ctrls_0_down_Decode_INSTRUCTION_0 = decode_ctrls_0_up_Decode_INSTRUCTION_0;
  assign decode_ctrls_0_down_Decode_DECOMPRESSION_FAULT_0 = decode_ctrls_0_up_Decode_DECOMPRESSION_FAULT_0;
  assign decode_ctrls_0_down_Decode_INSTRUCTION_RAW_0 = decode_ctrls_0_up_Decode_INSTRUCTION_RAW_0;
  assign decode_ctrls_0_down_Decode_INSTRUCTION_SLICE_COUNT_0 = decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0;
  assign decode_ctrls_0_down_PC_0 = decode_ctrls_0_up_PC_0;
  assign decode_ctrls_0_down_Decode_DOP_ID_0 = decode_ctrls_0_up_Decode_DOP_ID_0;
  assign decode_ctrls_0_down_Fetch_ID_0 = decode_ctrls_0_up_Fetch_ID_0;
  assign decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_0_0 = decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_0_0;
  assign decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_0_1 = decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_0_1;
  assign decode_ctrls_0_down_Prediction_BRANCH_HISTORY_0 = decode_ctrls_0_up_Prediction_BRANCH_HISTORY_0;
  assign decode_ctrls_0_down_TRAP_0 = decode_ctrls_0_up_TRAP_0;
  assign decode_ctrls_0_down_Prediction_ALIGNED_JUMPED_0 = decode_ctrls_0_up_Prediction_ALIGNED_JUMPED_0;
  assign decode_ctrls_0_down_Prediction_ALIGNED_JUMPED_PC_0 = decode_ctrls_0_up_Prediction_ALIGNED_JUMPED_PC_0;
  assign decode_ctrls_0_down_Prediction_ALIGNED_SLICES_BRANCH_0 = decode_ctrls_0_up_Prediction_ALIGNED_SLICES_BRANCH_0;
  assign decode_ctrls_0_down_Prediction_ALIGNED_SLICES_TAKEN_0 = decode_ctrls_0_up_Prediction_ALIGNED_SLICES_TAKEN_0;
  assign decode_ctrls_0_down_Prediction_ALIGN_REDO_0 = decode_ctrls_0_up_Prediction_ALIGN_REDO_0;
  assign decode_ctrls_1_down_valid = decode_ctrls_1_up_valid;
  assign decode_ctrls_1_up_ready = decode_ctrls_1_down_isReady;
  assign decode_ctrls_1_down_Decode_INSTRUCTION_0 = decode_ctrls_1_up_Decode_INSTRUCTION_0;
  assign decode_ctrls_1_down_Decode_DECOMPRESSION_FAULT_0 = decode_ctrls_1_up_Decode_DECOMPRESSION_FAULT_0;
  assign decode_ctrls_1_down_Decode_INSTRUCTION_RAW_0 = decode_ctrls_1_up_Decode_INSTRUCTION_RAW_0;
  assign decode_ctrls_1_down_Decode_INSTRUCTION_SLICE_COUNT_0 = decode_ctrls_1_up_Decode_INSTRUCTION_SLICE_COUNT_0;
  assign decode_ctrls_1_down_PC_0 = decode_ctrls_1_up_PC_0;
  assign decode_ctrls_1_down_Decode_DOP_ID_0 = decode_ctrls_1_up_Decode_DOP_ID_0;
  assign decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0_0 = decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_0_0;
  assign decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0_1 = decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_0_1;
  assign decode_ctrls_1_down_Prediction_BRANCH_HISTORY_0 = decode_ctrls_1_up_Prediction_BRANCH_HISTORY_0;
  assign decode_ctrls_1_down_Prediction_ALIGNED_JUMPED_0 = decode_ctrls_1_up_Prediction_ALIGNED_JUMPED_0;
  assign decode_ctrls_1_down_Prediction_ALIGNED_JUMPED_PC_0 = decode_ctrls_1_up_Prediction_ALIGNED_JUMPED_PC_0;
  assign decode_ctrls_1_down_Prediction_ALIGNED_SLICES_BRANCH_0 = decode_ctrls_1_up_Prediction_ALIGNED_SLICES_BRANCH_0;
  assign decode_ctrls_1_down_Prediction_ALIGNED_SLICES_TAKEN_0 = decode_ctrls_1_up_Prediction_ALIGNED_SLICES_TAKEN_0;
  assign decode_ctrls_1_down_Prediction_ALIGN_REDO_0 = decode_ctrls_1_up_Prediction_ALIGN_REDO_0;
  assign execute_ctrl0_down_ready = execute_ctrl1_up_ready;
  assign execute_ctrl1_down_ready = execute_ctrl2_up_ready;
  assign execute_ctrl2_down_ready = execute_ctrl3_up_ready;
  assign execute_ctrl3_down_ready = execute_ctrl4_up_ready;
  assign execute_ctrl4_down_ready = execute_ctrl5_up_ready;
  assign execute_ctrl0_up_ready = execute_ctrl0_down_isReady;
  assign execute_ctrl0_down_Decode_UOP_lane0 = execute_ctrl0_up_Decode_UOP_lane0;
  assign execute_ctrl0_down_Prediction_ALIGNED_JUMPED_lane0 = execute_ctrl0_up_Prediction_ALIGNED_JUMPED_lane0;
  assign execute_ctrl0_down_Prediction_ALIGNED_JUMPED_PC_lane0 = execute_ctrl0_up_Prediction_ALIGNED_JUMPED_PC_lane0;
  assign execute_ctrl0_down_Prediction_ALIGNED_SLICES_TAKEN_lane0 = execute_ctrl0_up_Prediction_ALIGNED_SLICES_TAKEN_lane0;
  assign execute_ctrl0_down_Prediction_ALIGNED_SLICES_BRANCH_lane0 = execute_ctrl0_up_Prediction_ALIGNED_SLICES_BRANCH_lane0;
  assign execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane0_0 = execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0;
  assign execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane0_1 = execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_1;
  assign execute_ctrl0_down_Prediction_BRANCH_HISTORY_lane0 = execute_ctrl0_up_Prediction_BRANCH_HISTORY_lane0;
  assign execute_ctrl0_down_Decode_INSTRUCTION_SLICE_COUNT_lane0 = execute_ctrl0_up_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  assign execute_ctrl0_down_PC_lane0 = execute_ctrl0_up_PC_lane0;
  assign execute_ctrl0_down_TRAP_lane0 = execute_ctrl0_up_TRAP_lane0;
  assign execute_ctrl0_down_Decode_UOP_ID_lane0 = execute_ctrl0_up_Decode_UOP_ID_lane0;
  assign execute_ctrl0_down_RS1_PHYS_lane0 = execute_ctrl0_up_RS1_PHYS_lane0;
  assign execute_ctrl0_down_RS2_PHYS_lane0 = execute_ctrl0_up_RS2_PHYS_lane0;
  assign execute_ctrl0_down_RD_PHYS_lane0 = execute_ctrl0_up_RD_PHYS_lane0;
  assign execute_ctrl0_down_COMPLETED_lane0 = execute_ctrl0_up_COMPLETED_lane0;
  assign execute_ctrl1_up_ready = execute_ctrl1_down_isReady;
  assign execute_ctrl1_down_Decode_UOP_lane0 = execute_ctrl1_up_Decode_UOP_lane0;
  assign execute_ctrl1_down_Prediction_ALIGNED_JUMPED_lane0 = execute_ctrl1_up_Prediction_ALIGNED_JUMPED_lane0;
  assign execute_ctrl1_down_Prediction_ALIGNED_JUMPED_PC_lane0 = execute_ctrl1_up_Prediction_ALIGNED_JUMPED_PC_lane0;
  assign execute_ctrl1_down_Prediction_ALIGNED_SLICES_TAKEN_lane0 = execute_ctrl1_up_Prediction_ALIGNED_SLICES_TAKEN_lane0;
  assign execute_ctrl1_down_Prediction_ALIGNED_SLICES_BRANCH_lane0 = execute_ctrl1_up_Prediction_ALIGNED_SLICES_BRANCH_lane0;
  assign execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane0_0 = execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane0_0;
  assign execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane0_1 = execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane0_1;
  assign execute_ctrl1_down_Prediction_BRANCH_HISTORY_lane0 = execute_ctrl1_up_Prediction_BRANCH_HISTORY_lane0;
  assign execute_ctrl1_down_Decode_INSTRUCTION_SLICE_COUNT_lane0 = execute_ctrl1_up_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  assign execute_ctrl1_down_PC_lane0 = execute_ctrl1_up_PC_lane0;
  assign execute_ctrl1_down_TRAP_lane0 = execute_ctrl1_up_TRAP_lane0;
  assign execute_ctrl1_down_Decode_UOP_ID_lane0 = execute_ctrl1_up_Decode_UOP_ID_lane0;
  assign execute_ctrl1_down_RS1_PHYS_lane0 = execute_ctrl1_up_RS1_PHYS_lane0;
  assign execute_ctrl1_down_RS2_PHYS_lane0 = execute_ctrl1_up_RS2_PHYS_lane0;
  assign execute_ctrl1_down_RD_PHYS_lane0 = execute_ctrl1_up_RD_PHYS_lane0;
  assign execute_ctrl1_down_COMPLETED_lane0 = execute_ctrl1_up_COMPLETED_lane0;
  assign execute_ctrl1_down_AguPlugin_SIZE_lane0 = execute_ctrl1_up_AguPlugin_SIZE_lane0;
  assign execute_ctrl2_up_ready = execute_ctrl2_down_isReady;
  assign execute_ctrl2_down_Decode_UOP_lane0 = execute_ctrl2_up_Decode_UOP_lane0;
  assign execute_ctrl2_down_Prediction_ALIGNED_JUMPED_lane0 = execute_ctrl2_up_Prediction_ALIGNED_JUMPED_lane0;
  assign execute_ctrl2_down_Prediction_ALIGNED_JUMPED_PC_lane0 = execute_ctrl2_up_Prediction_ALIGNED_JUMPED_PC_lane0;
  assign execute_ctrl2_down_Prediction_ALIGNED_SLICES_TAKEN_lane0 = execute_ctrl2_up_Prediction_ALIGNED_SLICES_TAKEN_lane0;
  assign execute_ctrl2_down_Prediction_ALIGNED_SLICES_BRANCH_lane0 = execute_ctrl2_up_Prediction_ALIGNED_SLICES_BRANCH_lane0;
  assign execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane0_0 = execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane0_0;
  assign execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane0_1 = execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane0_1;
  assign execute_ctrl2_down_Prediction_BRANCH_HISTORY_lane0 = execute_ctrl2_up_Prediction_BRANCH_HISTORY_lane0;
  assign execute_ctrl2_down_Decode_INSTRUCTION_SLICE_COUNT_lane0 = execute_ctrl2_up_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  assign execute_ctrl2_down_PC_lane0 = execute_ctrl2_up_PC_lane0;
  assign execute_ctrl2_down_Decode_UOP_ID_lane0 = execute_ctrl2_up_Decode_UOP_ID_lane0;
  assign execute_ctrl2_down_RD_PHYS_lane0 = execute_ctrl2_up_RD_PHYS_lane0;
  assign execute_ctrl2_down_AguPlugin_SIZE_lane0 = execute_ctrl2_up_AguPlugin_SIZE_lane0;
  assign execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0 = execute_ctrl2_up_early0_SrcPlugin_SRC1_lane0;
  assign execute_ctrl2_down_early0_SrcPlugin_SRC2_lane0 = execute_ctrl2_up_early0_SrcPlugin_SRC2_lane0;
  assign execute_ctrl2_down_integer_RS2_lane0 = execute_ctrl2_up_integer_RS2_lane0;
  assign execute_ctrl2_down_MAY_FLUSH_PRECISE_3_lane0 = execute_ctrl2_up_MAY_FLUSH_PRECISE_3_lane0;
  assign execute_ctrl2_down_early0_IntAluPlugin_SEL_lane0 = execute_ctrl2_up_early0_IntAluPlugin_SEL_lane0;
  assign execute_ctrl2_down_early0_BarrelShifterPlugin_SEL_lane0 = execute_ctrl2_up_early0_BarrelShifterPlugin_SEL_lane0;
  assign execute_ctrl2_down_early0_BranchPlugin_SEL_lane0 = execute_ctrl2_up_early0_BranchPlugin_SEL_lane0;
  assign execute_ctrl2_down_early0_MulPlugin_SEL_lane0 = execute_ctrl2_up_early0_MulPlugin_SEL_lane0;
  assign execute_ctrl2_down_early0_DivPlugin_SEL_lane0 = execute_ctrl2_up_early0_DivPlugin_SEL_lane0;
  assign execute_ctrl2_down_early0_EnvPlugin_SEL_lane0 = execute_ctrl2_up_early0_EnvPlugin_SEL_lane0;
  assign execute_ctrl2_down_MulPlugin_HIGH_lane0 = execute_ctrl2_up_MulPlugin_HIGH_lane0;
  assign execute_ctrl2_down_CsrAccessPlugin_SEL_lane0 = execute_ctrl2_up_CsrAccessPlugin_SEL_lane0;
  assign execute_ctrl2_down_AguPlugin_SEL_lane0 = execute_ctrl2_up_AguPlugin_SEL_lane0;
  assign execute_ctrl2_down_lane0_integer_WriteBackPlugin_SEL_lane0 = execute_ctrl2_up_lane0_integer_WriteBackPlugin_SEL_lane0;
  assign execute_ctrl2_down_COMPLETION_AT_2_lane0 = execute_ctrl2_up_COMPLETION_AT_2_lane0;
  assign execute_ctrl2_down_COMPLETION_AT_4_lane0 = execute_ctrl2_up_COMPLETION_AT_4_lane0;
  assign execute_ctrl2_down_COMPLETION_AT_3_lane0 = execute_ctrl2_up_COMPLETION_AT_3_lane0;
  assign execute_ctrl2_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0 = execute_ctrl2_up_lane0_logic_completions_onCtrl_0_ENABLE_lane0;
  assign execute_ctrl2_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0 = execute_ctrl2_up_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  assign execute_ctrl2_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0 = execute_ctrl2_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  assign execute_ctrl2_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0 = execute_ctrl2_up_early0_IntAluPlugin_ALU_ADD_SUB_lane0;
  assign execute_ctrl2_down_early0_IntAluPlugin_ALU_SLTX_lane0 = execute_ctrl2_up_early0_IntAluPlugin_ALU_SLTX_lane0;
  assign execute_ctrl2_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0 = execute_ctrl2_up_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  assign execute_ctrl2_down_SrcStageables_REVERT_lane0 = execute_ctrl2_up_SrcStageables_REVERT_lane0;
  assign execute_ctrl2_down_SrcStageables_ZERO_lane0 = execute_ctrl2_up_SrcStageables_ZERO_lane0;
  assign execute_ctrl2_down_lane0_IntFormatPlugin_logic_SIGNED_lane0 = execute_ctrl2_up_lane0_IntFormatPlugin_logic_SIGNED_lane0;
  assign execute_ctrl2_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0 = execute_ctrl2_up_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
  assign execute_ctrl2_down_BYPASSED_AT_3_lane0 = execute_ctrl2_up_BYPASSED_AT_3_lane0;
  assign execute_ctrl2_down_SrcStageables_UNSIGNED_lane0 = execute_ctrl2_up_SrcStageables_UNSIGNED_lane0;
  assign execute_ctrl2_down_BarrelShifterPlugin_LEFT_lane0 = execute_ctrl2_up_BarrelShifterPlugin_LEFT_lane0;
  assign execute_ctrl2_down_BarrelShifterPlugin_SIGNED_lane0 = execute_ctrl2_up_BarrelShifterPlugin_SIGNED_lane0;
  assign execute_ctrl2_down_BarrelShifterPlugin_IS_W_lane0 = execute_ctrl2_up_BarrelShifterPlugin_IS_W_lane0;
  assign execute_ctrl2_down_BarrelShifterPlugin_IS_W_RIGHT_lane0 = execute_ctrl2_up_BarrelShifterPlugin_IS_W_RIGHT_lane0;
  assign execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0 = execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane0;
  assign execute_ctrl2_down_RsUnsignedPlugin_RS1_SIGNED_lane0 = execute_ctrl2_up_RsUnsignedPlugin_RS1_SIGNED_lane0;
  assign execute_ctrl2_down_RsUnsignedPlugin_RS2_SIGNED_lane0 = execute_ctrl2_up_RsUnsignedPlugin_RS2_SIGNED_lane0;
  assign execute_ctrl2_down_DivPlugin_REM_lane0 = execute_ctrl2_up_DivPlugin_REM_lane0;
  assign execute_ctrl2_down_RsUnsignedPlugin_IS_W_lane0 = execute_ctrl2_up_RsUnsignedPlugin_IS_W_lane0;
  assign execute_ctrl2_down_CsrAccessPlugin_CSR_IMM_lane0 = execute_ctrl2_up_CsrAccessPlugin_CSR_IMM_lane0;
  assign execute_ctrl2_down_CsrAccessPlugin_CSR_MASK_lane0 = execute_ctrl2_up_CsrAccessPlugin_CSR_MASK_lane0;
  assign execute_ctrl2_down_CsrAccessPlugin_CSR_CLEAR_lane0 = execute_ctrl2_up_CsrAccessPlugin_CSR_CLEAR_lane0;
  assign execute_ctrl2_down_AguPlugin_LOAD_lane0 = execute_ctrl2_up_AguPlugin_LOAD_lane0;
  assign execute_ctrl2_down_AguPlugin_STORE_lane0 = execute_ctrl2_up_AguPlugin_STORE_lane0;
  assign execute_ctrl2_down_AguPlugin_ATOMIC_lane0 = execute_ctrl2_up_AguPlugin_ATOMIC_lane0;
  assign execute_ctrl2_down_AguPlugin_FLOAT_lane0 = execute_ctrl2_up_AguPlugin_FLOAT_lane0;
  assign execute_ctrl2_down_AguPlugin_CLEAN_lane0 = execute_ctrl2_up_AguPlugin_CLEAN_lane0;
  assign execute_ctrl2_down_AguPlugin_INVALIDATE_lane0 = execute_ctrl2_up_AguPlugin_INVALIDATE_lane0;
  assign execute_ctrl2_down_LsuPlugin_logic_LSU_PREFETCH_lane0 = execute_ctrl2_up_LsuPlugin_logic_LSU_PREFETCH_lane0;
  assign execute_ctrl2_down_early0_EnvPlugin_OP_lane0 = execute_ctrl2_up_early0_EnvPlugin_OP_lane0;
  assign execute_ctrl2_down_LsuL1Plugin_logic_FREEZE_HAZARD_lane0 = execute_ctrl2_up_LsuL1Plugin_logic_FREEZE_HAZARD_lane0;
  assign execute_ctrl3_up_ready = execute_ctrl3_down_isReady;
  assign execute_ctrl3_down_Decode_UOP_lane0 = execute_ctrl3_up_Decode_UOP_lane0;
  assign execute_ctrl3_down_Prediction_BRANCH_HISTORY_lane0 = execute_ctrl3_up_Prediction_BRANCH_HISTORY_lane0;
  assign execute_ctrl3_down_Decode_INSTRUCTION_SLICE_COUNT_lane0 = execute_ctrl3_up_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  assign execute_ctrl3_down_PC_lane0 = execute_ctrl3_up_PC_lane0;
  assign execute_ctrl3_down_TRAP_lane0 = execute_ctrl3_up_TRAP_lane0;
  assign execute_ctrl3_down_Decode_UOP_ID_lane0 = execute_ctrl3_up_Decode_UOP_ID_lane0;
  assign execute_ctrl3_down_RD_PHYS_lane0 = execute_ctrl3_up_RD_PHYS_lane0;
  assign execute_ctrl3_down_AguPlugin_SIZE_lane0 = execute_ctrl3_up_AguPlugin_SIZE_lane0;
  assign execute_ctrl3_down_integer_RS2_lane0 = execute_ctrl3_up_integer_RS2_lane0;
  assign execute_ctrl3_down_early0_MulPlugin_SEL_lane0 = execute_ctrl3_up_early0_MulPlugin_SEL_lane0;
  assign execute_ctrl3_down_early0_DivPlugin_SEL_lane0 = execute_ctrl3_up_early0_DivPlugin_SEL_lane0;
  assign execute_ctrl3_down_MulPlugin_HIGH_lane0 = execute_ctrl3_up_MulPlugin_HIGH_lane0;
  assign execute_ctrl3_down_CsrAccessPlugin_SEL_lane0 = execute_ctrl3_up_CsrAccessPlugin_SEL_lane0;
  assign execute_ctrl3_down_AguPlugin_SEL_lane0 = execute_ctrl3_up_AguPlugin_SEL_lane0;
  assign execute_ctrl3_down_LsuPlugin_logic_FENCE_lane0 = execute_ctrl3_up_LsuPlugin_logic_FENCE_lane0;
  assign execute_ctrl3_down_lane0_integer_WriteBackPlugin_SEL_lane0 = execute_ctrl3_up_lane0_integer_WriteBackPlugin_SEL_lane0;
  assign execute_ctrl3_down_COMPLETION_AT_4_lane0 = execute_ctrl3_up_COMPLETION_AT_4_lane0;
  assign execute_ctrl3_down_COMPLETION_AT_3_lane0 = execute_ctrl3_up_COMPLETION_AT_3_lane0;
  assign execute_ctrl3_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0 = execute_ctrl3_up_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  assign execute_ctrl3_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0 = execute_ctrl3_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  assign execute_ctrl3_down_lane0_IntFormatPlugin_logic_SIGNED_lane0 = execute_ctrl3_up_lane0_IntFormatPlugin_logic_SIGNED_lane0;
  assign execute_ctrl3_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0 = execute_ctrl3_up_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
  assign execute_ctrl3_down_AguPlugin_LOAD_lane0 = execute_ctrl3_up_AguPlugin_LOAD_lane0;
  assign execute_ctrl3_down_AguPlugin_STORE_lane0 = execute_ctrl3_up_AguPlugin_STORE_lane0;
  assign execute_ctrl3_down_AguPlugin_ATOMIC_lane0 = execute_ctrl3_up_AguPlugin_ATOMIC_lane0;
  assign execute_ctrl3_down_AguPlugin_FLOAT_lane0 = execute_ctrl3_up_AguPlugin_FLOAT_lane0;
  assign execute_ctrl3_down_LsuPlugin_logic_LSU_PREFETCH_lane0 = execute_ctrl3_up_LsuPlugin_logic_LSU_PREFETCH_lane0;
  assign execute_ctrl3_down_COMMIT_lane0 = execute_ctrl3_up_COMMIT_lane0;
  assign execute_ctrl3_down_early0_SrcPlugin_ADD_SUB_lane0 = execute_ctrl3_up_early0_SrcPlugin_ADD_SUB_lane0;
  assign execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0 = execute_ctrl3_up_LsuL1_MIXED_ADDRESS_lane0;
  assign execute_ctrl3_down_LsuL1Plugin_logic_BANK_BUSY_lane0 = execute_ctrl3_up_LsuL1Plugin_logic_BANK_BUSY_lane0;
  assign execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_VALID_lane0 = execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_VALID_lane0;
  assign execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_ADDRESS_lane0 = execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_ADDRESS_lane0;
  assign execute_ctrl3_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALID_lane0 = execute_ctrl3_up_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALID_lane0;
  assign execute_ctrl3_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_plru_0 = execute_ctrl3_up_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_plru_0;
  assign execute_ctrl3_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_dirty = execute_ctrl3_up_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_dirty;
  assign execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0 = execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0;
  assign execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0 = execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0;
  assign execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_0_lane0 = execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_0_lane0;
  assign execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_1_lane0 = execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_1_lane0;
  assign execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_2_lane0 = execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_2_lane0;
  assign execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_3_lane0 = execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_3_lane0;
  assign execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_4_lane0 = execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_4_lane0;
  assign execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_5_lane0 = execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_5_lane0;
  assign execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_6_lane0 = execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_6_lane0;
  assign execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_7_lane0 = execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_7_lane0;
  assign execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_8_lane0 = execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_8_lane0;
  assign execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_9_lane0 = execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_9_lane0;
  assign execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_10_lane0 = execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_10_lane0;
  assign execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_11_lane0 = execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_11_lane0;
  assign execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_12_lane0 = execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_12_lane0;
  assign execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_13_lane0 = execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_13_lane0;
  assign execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_14_lane0 = execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_14_lane0;
  assign execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_15_lane0 = execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_15_lane0;
  assign execute_ctrl3_down_DivPlugin_DIV_RESULT_lane0 = execute_ctrl3_up_DivPlugin_DIV_RESULT_lane0;
  assign execute_ctrl3_down_LsuPlugin_logic_FORCE_PHYSICAL_lane0 = execute_ctrl3_up_LsuPlugin_logic_FORCE_PHYSICAL_lane0;
  assign execute_ctrl3_down_LsuPlugin_logic_FROM_ACCESS_lane0 = execute_ctrl3_up_LsuPlugin_logic_FROM_ACCESS_lane0;
  assign execute_ctrl3_down_LsuL1_MASK_lane0 = execute_ctrl3_up_LsuL1_MASK_lane0;
  assign execute_ctrl3_down_LsuL1_SIZE_lane0 = execute_ctrl3_up_LsuL1_SIZE_lane0;
  assign execute_ctrl3_down_LsuL1_LOAD_lane0 = execute_ctrl3_up_LsuL1_LOAD_lane0;
  assign execute_ctrl3_down_LsuL1_ATOMIC_lane0 = execute_ctrl3_up_LsuL1_ATOMIC_lane0;
  assign execute_ctrl3_down_LsuL1_STORE_lane0 = execute_ctrl3_up_LsuL1_STORE_lane0;
  assign execute_ctrl3_down_LsuL1_CLEAN_lane0 = execute_ctrl3_up_LsuL1_CLEAN_lane0;
  assign execute_ctrl3_down_LsuL1_INVALID_lane0 = execute_ctrl3_up_LsuL1_INVALID_lane0;
  assign execute_ctrl3_down_LsuL1_PREFETCH_lane0 = execute_ctrl3_up_LsuL1_PREFETCH_lane0;
  assign execute_ctrl3_down_LsuL1_FLUSH_lane0 = execute_ctrl3_up_LsuL1_FLUSH_lane0;
  assign execute_ctrl3_down_Decode_STORE_ID_lane0 = execute_ctrl3_up_Decode_STORE_ID_lane0;
  assign execute_ctrl3_down_LsuPlugin_logic_FROM_LSU_lane0 = execute_ctrl3_up_LsuPlugin_logic_FROM_LSU_lane0;
  assign execute_ctrl3_down_LsuPlugin_logic_FROM_PREFETCH_lane0 = execute_ctrl3_up_LsuPlugin_logic_FROM_PREFETCH_lane0;
  assign execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_0_PERM_OK_lane0 = execute_ctrl3_up_LsuPlugin_logic_pmpPort_logic_onEntries_0_PERM_OK_lane0;
  assign execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_1_PERM_OK_lane0 = execute_ctrl3_up_LsuPlugin_logic_pmpPort_logic_onEntries_1_PERM_OK_lane0;
  assign execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_2_PERM_OK_lane0 = execute_ctrl3_up_LsuPlugin_logic_pmpPort_logic_onEntries_2_PERM_OK_lane0;
  assign execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_3_PERM_OK_lane0 = execute_ctrl3_up_LsuPlugin_logic_pmpPort_logic_onEntries_3_PERM_OK_lane0;
  assign execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_NEED_HIT_lane0 = execute_ctrl3_up_LsuPlugin_logic_pmpPort_logic_NEED_HIT_lane0;
  assign execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_valid = execute_ctrl3_up_MMU_L0_ENTRIES_lane0_0_valid;
  assign execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_virtualAddress = execute_ctrl3_up_MMU_L0_ENTRIES_lane0_0_virtualAddress;
  assign execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_physicalAddress = execute_ctrl3_up_MMU_L0_ENTRIES_lane0_0_physicalAddress;
  assign execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_allowRead = execute_ctrl3_up_MMU_L0_ENTRIES_lane0_0_allowRead;
  assign execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_allowWrite = execute_ctrl3_up_MMU_L0_ENTRIES_lane0_0_allowWrite;
  assign execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_allowExecute = execute_ctrl3_up_MMU_L0_ENTRIES_lane0_0_allowExecute;
  assign execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_allowUser = execute_ctrl3_up_MMU_L0_ENTRIES_lane0_0_allowUser;
  assign execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_valid = execute_ctrl3_up_MMU_L0_ENTRIES_lane0_1_valid;
  assign execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_virtualAddress = execute_ctrl3_up_MMU_L0_ENTRIES_lane0_1_virtualAddress;
  assign execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_physicalAddress = execute_ctrl3_up_MMU_L0_ENTRIES_lane0_1_physicalAddress;
  assign execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_allowRead = execute_ctrl3_up_MMU_L0_ENTRIES_lane0_1_allowRead;
  assign execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_allowWrite = execute_ctrl3_up_MMU_L0_ENTRIES_lane0_1_allowWrite;
  assign execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_allowExecute = execute_ctrl3_up_MMU_L0_ENTRIES_lane0_1_allowExecute;
  assign execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_allowUser = execute_ctrl3_up_MMU_L0_ENTRIES_lane0_1_allowUser;
  assign execute_ctrl3_down_MMU_L0_ENTRIES_lane0_2_valid = execute_ctrl3_up_MMU_L0_ENTRIES_lane0_2_valid;
  assign execute_ctrl3_down_MMU_L0_ENTRIES_lane0_2_virtualAddress = execute_ctrl3_up_MMU_L0_ENTRIES_lane0_2_virtualAddress;
  assign execute_ctrl3_down_MMU_L0_ENTRIES_lane0_2_physicalAddress = execute_ctrl3_up_MMU_L0_ENTRIES_lane0_2_physicalAddress;
  assign execute_ctrl3_down_MMU_L0_ENTRIES_lane0_2_allowRead = execute_ctrl3_up_MMU_L0_ENTRIES_lane0_2_allowRead;
  assign execute_ctrl3_down_MMU_L0_ENTRIES_lane0_2_allowWrite = execute_ctrl3_up_MMU_L0_ENTRIES_lane0_2_allowWrite;
  assign execute_ctrl3_down_MMU_L0_ENTRIES_lane0_2_allowExecute = execute_ctrl3_up_MMU_L0_ENTRIES_lane0_2_allowExecute;
  assign execute_ctrl3_down_MMU_L0_ENTRIES_lane0_2_allowUser = execute_ctrl3_up_MMU_L0_ENTRIES_lane0_2_allowUser;
  assign execute_ctrl3_down_MMU_L0_HITS_PRE_VALID_lane0 = execute_ctrl3_up_MMU_L0_HITS_PRE_VALID_lane0;
  assign execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_valid = execute_ctrl3_up_MMU_L1_ENTRIES_lane0_0_valid;
  assign execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_virtualAddress = execute_ctrl3_up_MMU_L1_ENTRIES_lane0_0_virtualAddress;
  assign execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_physicalAddress = execute_ctrl3_up_MMU_L1_ENTRIES_lane0_0_physicalAddress;
  assign execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_allowRead = execute_ctrl3_up_MMU_L1_ENTRIES_lane0_0_allowRead;
  assign execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_allowWrite = execute_ctrl3_up_MMU_L1_ENTRIES_lane0_0_allowWrite;
  assign execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_allowExecute = execute_ctrl3_up_MMU_L1_ENTRIES_lane0_0_allowExecute;
  assign execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_allowUser = execute_ctrl3_up_MMU_L1_ENTRIES_lane0_0_allowUser;
  assign execute_ctrl3_down_MMU_L1_HITS_PRE_VALID_lane0 = execute_ctrl3_up_MMU_L1_HITS_PRE_VALID_lane0;
  assign execute_ctrl4_up_ready = execute_ctrl4_down_isReady;
  assign execute_ctrl4_down_Decode_UOP_lane0 = execute_ctrl4_up_Decode_UOP_lane0;
  assign execute_ctrl4_down_Prediction_BRANCH_HISTORY_lane0 = execute_ctrl4_up_Prediction_BRANCH_HISTORY_lane0;
  assign execute_ctrl4_down_Decode_INSTRUCTION_SLICE_COUNT_lane0 = execute_ctrl4_up_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  assign execute_ctrl4_down_PC_lane0 = execute_ctrl4_up_PC_lane0;
  assign execute_ctrl4_down_Decode_UOP_ID_lane0 = execute_ctrl4_up_Decode_UOP_ID_lane0;
  assign execute_ctrl4_down_RD_PHYS_lane0 = execute_ctrl4_up_RD_PHYS_lane0;
  assign execute_ctrl4_down_AguPlugin_SIZE_lane0 = execute_ctrl4_up_AguPlugin_SIZE_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_SEL_lane0 = execute_ctrl4_up_early0_MulPlugin_SEL_lane0;
  assign execute_ctrl4_down_MulPlugin_HIGH_lane0 = execute_ctrl4_up_MulPlugin_HIGH_lane0;
  assign execute_ctrl4_down_AguPlugin_SEL_lane0 = execute_ctrl4_up_AguPlugin_SEL_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_FENCE_lane0 = execute_ctrl4_up_LsuPlugin_logic_FENCE_lane0;
  assign execute_ctrl4_down_lane0_integer_WriteBackPlugin_SEL_lane0 = execute_ctrl4_up_lane0_integer_WriteBackPlugin_SEL_lane0;
  assign execute_ctrl4_down_COMPLETION_AT_4_lane0 = execute_ctrl4_up_COMPLETION_AT_4_lane0;
  assign execute_ctrl4_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0 = execute_ctrl4_up_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  assign execute_ctrl4_down_lane0_IntFormatPlugin_logic_SIGNED_lane0 = execute_ctrl4_up_lane0_IntFormatPlugin_logic_SIGNED_lane0;
  assign execute_ctrl4_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0 = execute_ctrl4_up_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
  assign execute_ctrl4_down_AguPlugin_LOAD_lane0 = execute_ctrl4_up_AguPlugin_LOAD_lane0;
  assign execute_ctrl4_down_AguPlugin_STORE_lane0 = execute_ctrl4_up_AguPlugin_STORE_lane0;
  assign execute_ctrl4_down_AguPlugin_ATOMIC_lane0 = execute_ctrl4_up_AguPlugin_ATOMIC_lane0;
  assign execute_ctrl4_down_AguPlugin_FLOAT_lane0 = execute_ctrl4_up_AguPlugin_FLOAT_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_LSU_PREFETCH_lane0 = execute_ctrl4_up_LsuPlugin_logic_LSU_PREFETCH_lane0;
  assign execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0 = execute_ctrl4_up_LsuL1_MIXED_ADDRESS_lane0;
  assign execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0 = execute_ctrl4_up_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0;
  assign execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0 = execute_ctrl4_up_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_0_lane0 = execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_0_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_1_lane0 = execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_1_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_2_lane0 = execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_2_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_3_lane0 = execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_3_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_4_lane0 = execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_4_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_5_lane0 = execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_5_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_6_lane0 = execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_6_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_7_lane0 = execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_7_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_8_lane0 = execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_8_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_9_lane0 = execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_9_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_10_lane0 = execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_10_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_11_lane0 = execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_11_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_12_lane0 = execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_12_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_13_lane0 = execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_13_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_14_lane0 = execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_14_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_15_lane0 = execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_15_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_FROM_ACCESS_lane0 = execute_ctrl4_up_LsuPlugin_logic_FROM_ACCESS_lane0;
  assign execute_ctrl4_down_LsuL1_MASK_lane0 = execute_ctrl4_up_LsuL1_MASK_lane0;
  assign execute_ctrl4_down_LsuL1_SIZE_lane0 = execute_ctrl4_up_LsuL1_SIZE_lane0;
  assign execute_ctrl4_down_LsuL1_LOAD_lane0 = execute_ctrl4_up_LsuL1_LOAD_lane0;
  assign execute_ctrl4_down_LsuL1_ATOMIC_lane0 = execute_ctrl4_up_LsuL1_ATOMIC_lane0;
  assign execute_ctrl4_down_LsuL1_STORE_lane0 = execute_ctrl4_up_LsuL1_STORE_lane0;
  assign execute_ctrl4_down_LsuL1_CLEAN_lane0 = execute_ctrl4_up_LsuL1_CLEAN_lane0;
  assign execute_ctrl4_down_LsuL1_INVALID_lane0 = execute_ctrl4_up_LsuL1_INVALID_lane0;
  assign execute_ctrl4_down_LsuL1_PREFETCH_lane0 = execute_ctrl4_up_LsuL1_PREFETCH_lane0;
  assign execute_ctrl4_down_LsuL1_FLUSH_lane0 = execute_ctrl4_up_LsuL1_FLUSH_lane0;
  assign execute_ctrl4_down_Decode_STORE_ID_lane0 = execute_ctrl4_up_Decode_STORE_ID_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_FROM_LSU_lane0 = execute_ctrl4_up_LsuPlugin_logic_FROM_LSU_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_FROM_PREFETCH_lane0 = execute_ctrl4_up_LsuPlugin_logic_FROM_PREFETCH_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_0_PERM_OK_lane0 = execute_ctrl4_up_LsuPlugin_logic_pmpPort_logic_onEntries_0_PERM_OK_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_1_PERM_OK_lane0 = execute_ctrl4_up_LsuPlugin_logic_pmpPort_logic_onEntries_1_PERM_OK_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_2_PERM_OK_lane0 = execute_ctrl4_up_LsuPlugin_logic_pmpPort_logic_onEntries_2_PERM_OK_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_3_PERM_OK_lane0 = execute_ctrl4_up_LsuPlugin_logic_pmpPort_logic_onEntries_3_PERM_OK_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_NEED_HIT_lane0 = execute_ctrl4_up_LsuPlugin_logic_pmpPort_logic_NEED_HIT_lane0;
  assign execute_ctrl4_down_LsuL1Plugin_logic_SHARED_lane0_plru_0 = execute_ctrl4_up_LsuL1Plugin_logic_SHARED_lane0_plru_0;
  assign execute_ctrl4_down_LsuL1Plugin_logic_SHARED_lane0_dirty = execute_ctrl4_up_LsuL1Plugin_logic_SHARED_lane0_dirty;
  assign execute_ctrl4_down_LsuL1Plugin_logic_BANK_BUSY_REMAPPED_lane0 = execute_ctrl4_up_LsuL1Plugin_logic_BANK_BUSY_REMAPPED_lane0;
  assign execute_ctrl4_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0 = execute_ctrl4_up_LsuL1Plugin_logic_BANKS_MUXES_lane0_0;
  assign execute_ctrl4_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1 = execute_ctrl4_up_LsuL1Plugin_logic_BANKS_MUXES_lane0_1;
  assign execute_ctrl4_down_LsuL1Plugin_logic_WRITE_TO_READ_HAZARDS_lane0 = execute_ctrl4_up_LsuL1Plugin_logic_WRITE_TO_READ_HAZARDS_lane0;
  assign execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0 = execute_ctrl4_up_LsuL1_PHYSICAL_ADDRESS_lane0;
  assign execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_loaded = execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_loaded;
  assign execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_address = execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_address;
  assign execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault = execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault;
  assign execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_loaded = execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_loaded;
  assign execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_address = execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_address;
  assign execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault = execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault;
  assign execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0 = execute_ctrl4_up_LsuL1Plugin_logic_WAYS_HITS_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_logic_steps_0_adders_0_lane0 = execute_ctrl4_up_early0_MulPlugin_logic_steps_0_adders_0_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_logic_steps_0_adders_1_lane0 = execute_ctrl4_up_early0_MulPlugin_logic_steps_0_adders_1_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_logic_steps_0_adders_2_lane0 = execute_ctrl4_up_early0_MulPlugin_logic_steps_0_adders_2_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_onTrigger_HIT_lane0 = execute_ctrl4_up_LsuPlugin_logic_onTrigger_HIT_lane0;
  assign execute_ctrl4_down_MMU_TRANSLATED_lane0 = execute_ctrl4_up_MMU_TRANSLATED_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0 = execute_ctrl4_up_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_preCtrl_IS_AMO_lane0 = execute_ctrl4_up_LsuPlugin_logic_preCtrl_IS_AMO_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault = execute_ctrl4_up_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault;
  assign execute_ctrl4_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_io = execute_ctrl4_up_LsuPlugin_logic_onPma_CACHED_RSP_lane0_io;
  assign execute_ctrl4_down_LsuPlugin_logic_onPma_IO_RSP_lane0_fault = execute_ctrl4_up_LsuPlugin_logic_onPma_IO_RSP_lane0_fault;
  assign execute_ctrl4_down_LsuPlugin_logic_onPma_IO_RSP_lane0_io = execute_ctrl4_up_LsuPlugin_logic_onPma_IO_RSP_lane0_io;
  assign execute_ctrl4_down_LsuPlugin_logic_onPma_IO_lane0 = execute_ctrl4_up_LsuPlugin_logic_onPma_IO_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0 = execute_ctrl4_up_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_MMU_PAGE_FAULT_lane0 = execute_ctrl4_up_LsuPlugin_logic_MMU_PAGE_FAULT_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_MMU_FAILURE_lane0 = execute_ctrl4_up_LsuPlugin_logic_MMU_FAILURE_lane0;
  assign execute_ctrl4_down_MMU_ACCESS_FAULT_lane0 = execute_ctrl4_up_MMU_ACCESS_FAULT_lane0;
  assign execute_ctrl4_down_MMU_REFILL_lane0 = execute_ctrl4_up_MMU_REFILL_lane0;
  assign execute_ctrl4_down_MMU_HAZARD_lane0 = execute_ctrl4_up_MMU_HAZARD_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_0_napot_HIT_lane0 = execute_ctrl4_up_LsuPlugin_logic_pmpPort_logic_onEntries_0_napot_HIT_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_0_tor_BIGGER_lane0 = execute_ctrl4_up_LsuPlugin_logic_pmpPort_logic_onEntries_0_tor_BIGGER_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_1_napot_HIT_lane0 = execute_ctrl4_up_LsuPlugin_logic_pmpPort_logic_onEntries_1_napot_HIT_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_1_tor_BIGGER_lane0 = execute_ctrl4_up_LsuPlugin_logic_pmpPort_logic_onEntries_1_tor_BIGGER_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_2_napot_HIT_lane0 = execute_ctrl4_up_LsuPlugin_logic_pmpPort_logic_onEntries_2_napot_HIT_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_2_tor_BIGGER_lane0 = execute_ctrl4_up_LsuPlugin_logic_pmpPort_logic_onEntries_2_tor_BIGGER_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_3_napot_HIT_lane0 = execute_ctrl4_up_LsuPlugin_logic_pmpPort_logic_onEntries_3_napot_HIT_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_pmpPort_logic_onEntries_3_tor_BIGGER_lane0 = execute_ctrl4_up_LsuPlugin_logic_pmpPort_logic_onEntries_3_tor_BIGGER_lane0;
  assign execute_ctrl4_down_MMU_BYPASS_TRANSLATION_lane0 = execute_ctrl4_up_MMU_BYPASS_TRANSLATION_lane0;
  assign execute_ctrl5_up_ready = execute_ctrl5_down_isReady;
  assign execute_ctrl5_down_LANE_SEL_lane0 = execute_ctrl5_up_LANE_SEL_lane0;
  assign execute_ctrl5_down_RD_PHYS_lane0 = execute_ctrl5_up_RD_PHYS_lane0;
  assign execute_ctrl5_down_COMMIT_lane0 = execute_ctrl5_up_COMMIT_lane0;
  assign execute_ctrl5_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 = execute_ctrl5_up_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
  assign fetch_logic_ctrls_0_down_isFiring = (fetch_logic_ctrls_0_down_isValid && fetch_logic_ctrls_0_down_isReady);
  assign fetch_logic_ctrls_0_down_isValid = fetch_logic_ctrls_0_down_valid;
  assign fetch_logic_ctrls_0_down_isReady = fetch_logic_ctrls_0_down_ready;
  assign fetch_logic_ctrls_1_up_isValid = fetch_logic_ctrls_1_up_valid;
  assign fetch_logic_ctrls_1_up_isReady = fetch_logic_ctrls_1_up_ready;
  assign fetch_logic_ctrls_1_up_isCancel = fetch_logic_ctrls_1_up_cancel;
  assign fetch_logic_ctrls_1_down_isValid = fetch_logic_ctrls_1_down_valid;
  assign fetch_logic_ctrls_1_down_isReady = fetch_logic_ctrls_1_down_ready;
  assign fetch_logic_ctrls_2_up_isMoving = (fetch_logic_ctrls_2_up_isValid && (fetch_logic_ctrls_2_up_isReady || fetch_logic_ctrls_2_up_isCancel));
  assign fetch_logic_ctrls_2_up_isValid = fetch_logic_ctrls_2_up_valid;
  assign fetch_logic_ctrls_2_up_isReady = fetch_logic_ctrls_2_up_ready;
  assign fetch_logic_ctrls_2_up_isCancel = fetch_logic_ctrls_2_up_cancel;
  assign fetch_logic_ctrls_2_up_isCanceling = (fetch_logic_ctrls_2_up_isValid && fetch_logic_ctrls_2_up_isCancel);
  assign fetch_logic_ctrls_0_up_isFiring = (fetch_logic_ctrls_0_up_isValid && fetch_logic_ctrls_0_up_isReady);
  assign fetch_logic_ctrls_0_up_isValid = fetch_logic_ctrls_0_up_valid;
  assign fetch_logic_ctrls_0_up_isReady = fetch_logic_ctrls_0_up_ready;
  assign fetch_logic_ctrls_2_down_isValid = fetch_logic_ctrls_2_down_valid;
  assign fetch_logic_ctrls_2_down_isReady = fetch_logic_ctrls_2_down_ready;
  assign fetch_logic_ctrls_2_down_isCancel = 1'b0;
  assign decode_ctrls_0_down_isValid = decode_ctrls_0_down_valid;
  assign decode_ctrls_0_down_isReady = decode_ctrls_0_down_ready;
  assign decode_ctrls_1_up_isMoving = (decode_ctrls_1_up_isValid && decode_ctrls_1_up_isReady);
  assign decode_ctrls_1_up_isValid = decode_ctrls_1_up_valid;
  assign decode_ctrls_1_up_isReady = decode_ctrls_1_up_ready;
  assign decode_ctrls_1_up_isCanceling = 1'b0;
  assign decode_ctrls_0_up_isFiring = (decode_ctrls_0_up_isValid && decode_ctrls_0_up_isReady);
  assign decode_ctrls_0_up_isMoving = (decode_ctrls_0_up_isValid && decode_ctrls_0_up_isReady);
  assign decode_ctrls_0_up_isValid = decode_ctrls_0_up_valid;
  assign decode_ctrls_0_up_isReady = decode_ctrls_0_up_ready;
  assign decode_ctrls_0_up_isCancel = 1'b0;
  assign decode_ctrls_1_down_isReady = decode_ctrls_1_down_ready;
  assign execute_ctrl0_down_isReady = execute_ctrl0_down_ready;
  assign execute_ctrl1_down_isReady = execute_ctrl1_down_ready;
  assign execute_ctrl2_down_isReady = execute_ctrl2_down_ready;
  assign execute_ctrl3_down_isReady = execute_ctrl3_down_ready;
  assign execute_ctrl4_up_isReady = execute_ctrl4_up_ready;
  assign execute_ctrl4_down_isReady = execute_ctrl4_down_ready;
  assign execute_ctrl5_down_isReady = execute_ctrl5_down_ready;
  always @(*) begin
    LsuPlugin_logic_flusher_stateNext = LsuPlugin_logic_flusher_stateReg;
    case(LsuPlugin_logic_flusher_stateReg)
      LsuPlugin_logic_flusher_CMD : begin
        if(when_LsuPlugin_l368) begin
          LsuPlugin_logic_flusher_stateNext = LsuPlugin_logic_flusher_COMPLETION;
        end
      end
      LsuPlugin_logic_flusher_COMPLETION : begin
        if(when_LsuPlugin_l376) begin
          LsuPlugin_logic_flusher_stateNext = LsuPlugin_logic_flusher_IDLE;
        end
      end
      default : begin
        if(LsuPlugin_logic_flusher_arbiter_io_output_valid) begin
          LsuPlugin_logic_flusher_stateNext = LsuPlugin_logic_flusher_CMD;
        end
      end
    endcase
    if(LsuPlugin_logic_flusher_wantKill) begin
      LsuPlugin_logic_flusher_stateNext = LsuPlugin_logic_flusher_IDLE;
    end
  end

  assign when_LsuPlugin_l368 = (LsuPlugin_logic_flusher_cmdCounter[6] && (! LsuPlugin_logic_flusher_inflight));
  assign when_LsuPlugin_l376 = (! (|LsuPlugin_logic_flusher_waiter));
  assign LsuPlugin_logic_flusher_onExit_IDLE = ((LsuPlugin_logic_flusher_stateNext != LsuPlugin_logic_flusher_IDLE) && (LsuPlugin_logic_flusher_stateReg == LsuPlugin_logic_flusher_IDLE));
  assign LsuPlugin_logic_flusher_onExit_CMD = ((LsuPlugin_logic_flusher_stateNext != LsuPlugin_logic_flusher_CMD) && (LsuPlugin_logic_flusher_stateReg == LsuPlugin_logic_flusher_CMD));
  assign LsuPlugin_logic_flusher_onExit_COMPLETION = ((LsuPlugin_logic_flusher_stateNext != LsuPlugin_logic_flusher_COMPLETION) && (LsuPlugin_logic_flusher_stateReg == LsuPlugin_logic_flusher_COMPLETION));
  assign LsuPlugin_logic_flusher_onEntry_IDLE = ((LsuPlugin_logic_flusher_stateNext == LsuPlugin_logic_flusher_IDLE) && (LsuPlugin_logic_flusher_stateReg != LsuPlugin_logic_flusher_IDLE));
  assign LsuPlugin_logic_flusher_onEntry_CMD = ((LsuPlugin_logic_flusher_stateNext == LsuPlugin_logic_flusher_CMD) && (LsuPlugin_logic_flusher_stateReg != LsuPlugin_logic_flusher_CMD));
  assign LsuPlugin_logic_flusher_onEntry_COMPLETION = ((LsuPlugin_logic_flusher_stateNext == LsuPlugin_logic_flusher_COMPLETION) && (LsuPlugin_logic_flusher_stateReg != LsuPlugin_logic_flusher_COMPLETION));
  always @(*) begin
    TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_stateReg;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
        if(TrapPlugin_logic_harts_0_trap_trigger_valid) begin
          TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_COMPUTE;
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
        if(when_TrapPlugin_l453) begin
          TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL;
        end else begin
          case(TrapPlugin_logic_harts_0_trap_pending_state_code)
            4'b0000 : begin
              TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_RUNNING;
            end
            4'b0001 : begin
              if(when_TrapPlugin_l481) begin
                TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC;
              end
            end
            4'b0010 : begin
              TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH;
            end
            4'b0100 : begin
              TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_JUMP;
            end
            4'b0101 : begin
              TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_JUMP;
            end
            4'b1000 : begin
              if(TrapPlugin_api_harts_0_askWake) begin
                TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_JUMP;
              end
            end
            4'b0110 : begin
              if(TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidate_cmd_ready) begin
                TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_JUMP;
              end
            end
            4'b0111 : begin
              if(TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_cmd_ready) begin
                TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP;
              end
            end
            default : begin
            end
          endcase
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
        if(TrapPlugin_logic_harts_0_crsPorts_write_ready) begin
          TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC;
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
        if(TrapPlugin_logic_harts_0_crsPorts_write_ready) begin
          TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC;
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
        if(TrapPlugin_logic_harts_0_crsPorts_read_ready) begin
          TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_TRAP_WAIT;
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_WAIT : begin
        if(when_TrapPlugin_l615) begin
          TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY;
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
        TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_RUNNING;
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
        if(TrapPlugin_logic_harts_0_crsPorts_read_ready) begin
          TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY;
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
        TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_RUNNING;
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
        if(TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_valid) begin
          TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_JUMP;
          if(when_TrapPlugin_l555) begin
            TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL;
          end
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
        TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_RUNNING;
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
        if(TrapPlugin_logic_lsuL1Invalidate_0_cmd_ready) begin
          TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH;
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
        if(TrapPlugin_logic_fetchL1Invalidate_0_cmd_ready) begin
          TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_JUMP;
        end
      end
      default : begin
        if(when_TrapPlugin_l406) begin
          TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_RUNNING;
        end
      end
    endcase
    if(TrapPlugin_logic_harts_0_trap_fsm_wantKill) begin
      TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_RESET;
    end
  end

  assign when_TrapPlugin_l453 = ((TrapPlugin_logic_harts_0_trap_pending_state_exception || TrapPlugin_logic_harts_0_trap_fsm_triggerEbreak) || TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_interrupt);
  assign when_TrapPlugin_l481 = (! TrapPlugin_api_harts_0_holdPrivChange);
  always @(*) begin
    _zz_TrapPlugin_logic_harts_0_crsPorts_write_address = 4'b0111;
    case(TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_targetPrivilege)
      2'b01 : begin
        _zz_TrapPlugin_logic_harts_0_crsPorts_write_address = 4'b0011;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_TrapPlugin_logic_harts_0_crsPorts_write_address_1 = 4'b1000;
    case(TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_targetPrivilege)
      2'b01 : begin
        _zz_TrapPlugin_logic_harts_0_crsPorts_write_address_1 = 4'b0100;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_TrapPlugin_logic_harts_0_crsPorts_read_address = 4'b1001;
    case(TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_targetPrivilege)
      2'b01 : begin
        _zz_TrapPlugin_logic_harts_0_crsPorts_read_address = 4'b0101;
      end
      default : begin
      end
    endcase
  end

  assign when_TrapPlugin_l615 = (! TrapPlugin_api_harts_0_holdPrivChange);
  always @(*) begin
    _zz_TrapPlugin_logic_harts_0_crsPorts_read_address_1 = 4'b0111;
    case(TrapPlugin_logic_harts_0_trap_fsm_xretPrivilege)
      2'b01 : begin
        _zz_TrapPlugin_logic_harts_0_crsPorts_read_address_1 = 4'b0011;
      end
      default : begin
      end
    endcase
  end

  assign when_TrapPlugin_l712 = (TrapPlugin_logic_harts_0_trap_pending_xret_targetPrivilege != 2'b11);
  assign switch_TrapPlugin_l713 = TrapPlugin_logic_harts_0_trap_pending_state_arg[1 : 0];
  assign when_TrapPlugin_l555 = (bits_pageFault || bits_accessFault);
  assign switch_TrapPlugin_l557 = {bits_accessFault,TrapPlugin_logic_harts_0_trap_pending_state_arg[1 : 0]};
  assign when_TrapPlugin_l406 = (&{TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidated,TrapPlugin_logic_harts_0_trap_fsm_resetToRunConditions_0});
  assign TrapPlugin_logic_harts_0_trap_fsm_onExit_RESET = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext != TrapPlugin_logic_harts_0_trap_fsm_RESET) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_RESET));
  assign TrapPlugin_logic_harts_0_trap_fsm_onExit_RUNNING = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext != TrapPlugin_logic_harts_0_trap_fsm_RUNNING) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_RUNNING));
  assign TrapPlugin_logic_harts_0_trap_fsm_onExit_COMPUTE = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext != TrapPlugin_logic_harts_0_trap_fsm_COMPUTE) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_COMPUTE));
  assign TrapPlugin_logic_harts_0_trap_fsm_onExit_TRAP_EPC = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext != TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC));
  assign TrapPlugin_logic_harts_0_trap_fsm_onExit_TRAP_TVAL = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext != TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL));
  assign TrapPlugin_logic_harts_0_trap_fsm_onExit_TRAP_TVEC = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext != TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC));
  assign TrapPlugin_logic_harts_0_trap_fsm_onExit_TRAP_WAIT = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext != TrapPlugin_logic_harts_0_trap_fsm_TRAP_WAIT) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_TRAP_WAIT));
  assign TrapPlugin_logic_harts_0_trap_fsm_onExit_TRAP_APPLY = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext != TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY));
  assign TrapPlugin_logic_harts_0_trap_fsm_onExit_XRET_EPC = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext != TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC));
  assign TrapPlugin_logic_harts_0_trap_fsm_onExit_XRET_APPLY = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext != TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY));
  assign TrapPlugin_logic_harts_0_trap_fsm_onExit_ATS_RSP = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext != TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP));
  assign TrapPlugin_logic_harts_0_trap_fsm_onExit_JUMP = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext != TrapPlugin_logic_harts_0_trap_fsm_JUMP) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_JUMP));
  assign TrapPlugin_logic_harts_0_trap_fsm_onExit_LSU_FLUSH = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext != TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH));
  assign TrapPlugin_logic_harts_0_trap_fsm_onExit_FETCH_FLUSH = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext != TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH));
  assign TrapPlugin_logic_harts_0_trap_fsm_onEntry_RESET = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext == TrapPlugin_logic_harts_0_trap_fsm_RESET) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg != TrapPlugin_logic_harts_0_trap_fsm_RESET));
  assign TrapPlugin_logic_harts_0_trap_fsm_onEntry_RUNNING = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext == TrapPlugin_logic_harts_0_trap_fsm_RUNNING) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg != TrapPlugin_logic_harts_0_trap_fsm_RUNNING));
  assign TrapPlugin_logic_harts_0_trap_fsm_onEntry_COMPUTE = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext == TrapPlugin_logic_harts_0_trap_fsm_COMPUTE) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg != TrapPlugin_logic_harts_0_trap_fsm_COMPUTE));
  assign TrapPlugin_logic_harts_0_trap_fsm_onEntry_TRAP_EPC = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext == TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg != TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC));
  assign TrapPlugin_logic_harts_0_trap_fsm_onEntry_TRAP_TVAL = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext == TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg != TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL));
  assign TrapPlugin_logic_harts_0_trap_fsm_onEntry_TRAP_TVEC = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext == TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg != TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC));
  assign TrapPlugin_logic_harts_0_trap_fsm_onEntry_TRAP_WAIT = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext == TrapPlugin_logic_harts_0_trap_fsm_TRAP_WAIT) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg != TrapPlugin_logic_harts_0_trap_fsm_TRAP_WAIT));
  assign TrapPlugin_logic_harts_0_trap_fsm_onEntry_TRAP_APPLY = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext == TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg != TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY));
  assign TrapPlugin_logic_harts_0_trap_fsm_onEntry_XRET_EPC = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext == TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg != TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC));
  assign TrapPlugin_logic_harts_0_trap_fsm_onEntry_XRET_APPLY = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext == TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg != TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY));
  assign TrapPlugin_logic_harts_0_trap_fsm_onEntry_ATS_RSP = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext == TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg != TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP));
  assign TrapPlugin_logic_harts_0_trap_fsm_onEntry_JUMP = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext == TrapPlugin_logic_harts_0_trap_fsm_JUMP) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg != TrapPlugin_logic_harts_0_trap_fsm_JUMP));
  assign TrapPlugin_logic_harts_0_trap_fsm_onEntry_LSU_FLUSH = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext == TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg != TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH));
  assign TrapPlugin_logic_harts_0_trap_fsm_onEntry_FETCH_FLUSH = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext == TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg != TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH));
  always @(*) begin
    MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_stateReg;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
        if(MmuPlugin_logic_refill_arbiter_io_output_valid) begin
          MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_CMD_2;
        end
      end
      MmuPlugin_logic_refill_CMD_0 : begin
        if(when_MmuPlugin_l516) begin
          if(MmuPlugin_logic_accessBus_cmd_ready) begin
            MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_RSP_0;
          end
        end
      end
      MmuPlugin_logic_refill_CMD_1 : begin
        if(when_MmuPlugin_l516_1) begin
          if(MmuPlugin_logic_accessBus_cmd_ready) begin
            MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_RSP_1;
          end
        end
      end
      MmuPlugin_logic_refill_CMD_2 : begin
        if(when_MmuPlugin_l516_2) begin
          if(MmuPlugin_logic_accessBus_cmd_ready) begin
            MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_RSP_2;
          end
        end
      end
      MmuPlugin_logic_refill_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_CMD_0;
          end else begin
            MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_DONE_0;
          end
        end
      end
      MmuPlugin_logic_refill_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_CMD_1;
          end else begin
            if(when_MmuPlugin_l534) begin
              MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_DONE_1;
            end else begin
              MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_CMD_0;
            end
          end
        end
      end
      MmuPlugin_logic_refill_RSP_2 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_CMD_2;
          end else begin
            if(when_MmuPlugin_l534_1) begin
              MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_DONE_2;
            end else begin
              MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_CMD_1;
            end
          end
        end
      end
      MmuPlugin_logic_refill_DONE_0 : begin
        MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_IDLE;
      end
      MmuPlugin_logic_refill_DONE_1 : begin
        MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_IDLE;
      end
      MmuPlugin_logic_refill_DONE_2 : begin
        MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_IDLE;
      end
      default : begin
      end
    endcase
    if(MmuPlugin_logic_refill_wantStart) begin
      MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_IDLE;
    end
    if(MmuPlugin_logic_refill_wantKill) begin
      MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_BOOT;
    end
  end

  assign when_MmuPlugin_l516 = (1'b1 && (MmuPlugin_logic_refill_cacheRefillAny == 1'b0));
  assign when_MmuPlugin_l516_1 = (1'b1 && (MmuPlugin_logic_refill_cacheRefillAny == 1'b0));
  assign when_MmuPlugin_l516_2 = (1'b1 && (MmuPlugin_logic_refill_cacheRefillAny == 1'b0));
  assign when_MmuPlugin_l525 = (! MmuPlugin_logic_refill_load_leaf);
  assign when_MmuPlugin_l534 = (MmuPlugin_logic_refill_load_leaf || MmuPlugin_logic_refill_load_exception);
  assign when_MmuPlugin_l534_1 = (MmuPlugin_logic_refill_load_leaf || MmuPlugin_logic_refill_load_exception);
  assign _zz_55 = MmuPlugin_logic_refill_portOhReg[0];
  assign when_MmuPlugin_l505 = ((MmuPlugin_logic_refill_fetch_0_pageFault || MmuPlugin_logic_refill_fetch_0_accessFault) || (! MmuPlugin_logic_refill_storageEnable));
  assign when_MmuPlugin_l505_1 = ((MmuPlugin_logic_refill_fetch_0_pageFault || MmuPlugin_logic_refill_fetch_0_accessFault) || (! MmuPlugin_logic_refill_storageEnable));
  assign when_MmuPlugin_l505_2 = ((MmuPlugin_logic_refill_fetch_1_pageFault || MmuPlugin_logic_refill_fetch_1_accessFault) || (! MmuPlugin_logic_refill_storageEnable));
  assign when_MmuPlugin_l505_3 = ((MmuPlugin_logic_refill_fetch_1_pageFault || MmuPlugin_logic_refill_fetch_1_accessFault) || (! MmuPlugin_logic_refill_storageEnable));
  assign when_MmuPlugin_l505_4 = ((MmuPlugin_logic_refill_fetch_2_pageFault || MmuPlugin_logic_refill_fetch_2_accessFault) || (! MmuPlugin_logic_refill_storageEnable));
  assign when_MmuPlugin_l505_5 = ((MmuPlugin_logic_refill_fetch_2_pageFault || MmuPlugin_logic_refill_fetch_2_accessFault) || (! MmuPlugin_logic_refill_storageEnable));
  assign MmuPlugin_logic_refill_onExit_BOOT = ((MmuPlugin_logic_refill_stateNext != MmuPlugin_logic_refill_BOOT) && (MmuPlugin_logic_refill_stateReg == MmuPlugin_logic_refill_BOOT));
  assign MmuPlugin_logic_refill_onExit_IDLE = ((MmuPlugin_logic_refill_stateNext != MmuPlugin_logic_refill_IDLE) && (MmuPlugin_logic_refill_stateReg == MmuPlugin_logic_refill_IDLE));
  assign MmuPlugin_logic_refill_onExit_CMD_0 = ((MmuPlugin_logic_refill_stateNext != MmuPlugin_logic_refill_CMD_0) && (MmuPlugin_logic_refill_stateReg == MmuPlugin_logic_refill_CMD_0));
  assign MmuPlugin_logic_refill_onExit_CMD_1 = ((MmuPlugin_logic_refill_stateNext != MmuPlugin_logic_refill_CMD_1) && (MmuPlugin_logic_refill_stateReg == MmuPlugin_logic_refill_CMD_1));
  assign MmuPlugin_logic_refill_onExit_CMD_2 = ((MmuPlugin_logic_refill_stateNext != MmuPlugin_logic_refill_CMD_2) && (MmuPlugin_logic_refill_stateReg == MmuPlugin_logic_refill_CMD_2));
  assign MmuPlugin_logic_refill_onExit_RSP_0 = ((MmuPlugin_logic_refill_stateNext != MmuPlugin_logic_refill_RSP_0) && (MmuPlugin_logic_refill_stateReg == MmuPlugin_logic_refill_RSP_0));
  assign MmuPlugin_logic_refill_onExit_RSP_1 = ((MmuPlugin_logic_refill_stateNext != MmuPlugin_logic_refill_RSP_1) && (MmuPlugin_logic_refill_stateReg == MmuPlugin_logic_refill_RSP_1));
  assign MmuPlugin_logic_refill_onExit_RSP_2 = ((MmuPlugin_logic_refill_stateNext != MmuPlugin_logic_refill_RSP_2) && (MmuPlugin_logic_refill_stateReg == MmuPlugin_logic_refill_RSP_2));
  assign MmuPlugin_logic_refill_onExit_DONE_0 = ((MmuPlugin_logic_refill_stateNext != MmuPlugin_logic_refill_DONE_0) && (MmuPlugin_logic_refill_stateReg == MmuPlugin_logic_refill_DONE_0));
  assign MmuPlugin_logic_refill_onExit_DONE_1 = ((MmuPlugin_logic_refill_stateNext != MmuPlugin_logic_refill_DONE_1) && (MmuPlugin_logic_refill_stateReg == MmuPlugin_logic_refill_DONE_1));
  assign MmuPlugin_logic_refill_onExit_DONE_2 = ((MmuPlugin_logic_refill_stateNext != MmuPlugin_logic_refill_DONE_2) && (MmuPlugin_logic_refill_stateReg == MmuPlugin_logic_refill_DONE_2));
  assign MmuPlugin_logic_refill_onEntry_BOOT = ((MmuPlugin_logic_refill_stateNext == MmuPlugin_logic_refill_BOOT) && (MmuPlugin_logic_refill_stateReg != MmuPlugin_logic_refill_BOOT));
  assign MmuPlugin_logic_refill_onEntry_IDLE = ((MmuPlugin_logic_refill_stateNext == MmuPlugin_logic_refill_IDLE) && (MmuPlugin_logic_refill_stateReg != MmuPlugin_logic_refill_IDLE));
  assign MmuPlugin_logic_refill_onEntry_CMD_0 = ((MmuPlugin_logic_refill_stateNext == MmuPlugin_logic_refill_CMD_0) && (MmuPlugin_logic_refill_stateReg != MmuPlugin_logic_refill_CMD_0));
  assign MmuPlugin_logic_refill_onEntry_CMD_1 = ((MmuPlugin_logic_refill_stateNext == MmuPlugin_logic_refill_CMD_1) && (MmuPlugin_logic_refill_stateReg != MmuPlugin_logic_refill_CMD_1));
  assign MmuPlugin_logic_refill_onEntry_CMD_2 = ((MmuPlugin_logic_refill_stateNext == MmuPlugin_logic_refill_CMD_2) && (MmuPlugin_logic_refill_stateReg != MmuPlugin_logic_refill_CMD_2));
  assign MmuPlugin_logic_refill_onEntry_RSP_0 = ((MmuPlugin_logic_refill_stateNext == MmuPlugin_logic_refill_RSP_0) && (MmuPlugin_logic_refill_stateReg != MmuPlugin_logic_refill_RSP_0));
  assign MmuPlugin_logic_refill_onEntry_RSP_1 = ((MmuPlugin_logic_refill_stateNext == MmuPlugin_logic_refill_RSP_1) && (MmuPlugin_logic_refill_stateReg != MmuPlugin_logic_refill_RSP_1));
  assign MmuPlugin_logic_refill_onEntry_RSP_2 = ((MmuPlugin_logic_refill_stateNext == MmuPlugin_logic_refill_RSP_2) && (MmuPlugin_logic_refill_stateReg != MmuPlugin_logic_refill_RSP_2));
  assign MmuPlugin_logic_refill_onEntry_DONE_0 = ((MmuPlugin_logic_refill_stateNext == MmuPlugin_logic_refill_DONE_0) && (MmuPlugin_logic_refill_stateReg != MmuPlugin_logic_refill_DONE_0));
  assign MmuPlugin_logic_refill_onEntry_DONE_1 = ((MmuPlugin_logic_refill_stateNext == MmuPlugin_logic_refill_DONE_1) && (MmuPlugin_logic_refill_stateReg != MmuPlugin_logic_refill_DONE_1));
  assign MmuPlugin_logic_refill_onEntry_DONE_2 = ((MmuPlugin_logic_refill_stateNext == MmuPlugin_logic_refill_DONE_2) && (MmuPlugin_logic_refill_stateReg != MmuPlugin_logic_refill_DONE_2));
  always @(*) begin
    PerformanceCounterPlugin_logic_fsm_stateNext = PerformanceCounterPlugin_logic_fsm_stateReg;
    case(PerformanceCounterPlugin_logic_fsm_stateReg)
      PerformanceCounterPlugin_logic_fsm_IDLE : begin
        if(PerformanceCounterPlugin_logic_fsm_csrWriteCmd_valid) begin
          PerformanceCounterPlugin_logic_fsm_stateNext = PerformanceCounterPlugin_logic_fsm_CSR_WRITE;
        end else begin
          if(PerformanceCounterPlugin_logic_fsm_flusherCmd_valid) begin
            PerformanceCounterPlugin_logic_fsm_stateNext = PerformanceCounterPlugin_logic_fsm_READ_LOW;
          end else begin
            if(PerformanceCounterPlugin_logic_fsm_csrReadCmd_valid) begin
              PerformanceCounterPlugin_logic_fsm_stateNext = PerformanceCounterPlugin_logic_fsm_READ_LOW;
            end
          end
        end
      end
      PerformanceCounterPlugin_logic_fsm_READ_LOW : begin
        if(PerformanceCounterPlugin_logic_readPort_ready) begin
          PerformanceCounterPlugin_logic_fsm_stateNext = PerformanceCounterPlugin_logic_fsm_CALC_LOW;
        end
      end
      PerformanceCounterPlugin_logic_fsm_CALC_LOW : begin
        if(PerformanceCounterPlugin_logic_writePort_ready) begin
          PerformanceCounterPlugin_logic_fsm_stateNext = PerformanceCounterPlugin_logic_fsm_IDLE;
        end
      end
      PerformanceCounterPlugin_logic_fsm_CSR_WRITE : begin
        PerformanceCounterPlugin_logic_fsm_stateNext = PerformanceCounterPlugin_logic_fsm_IDLE;
      end
      default : begin
      end
    endcase
    if(PerformanceCounterPlugin_logic_fsm_wantStart) begin
      PerformanceCounterPlugin_logic_fsm_stateNext = PerformanceCounterPlugin_logic_fsm_IDLE;
    end
    if(PerformanceCounterPlugin_logic_fsm_wantKill) begin
      PerformanceCounterPlugin_logic_fsm_stateNext = PerformanceCounterPlugin_logic_fsm_BOOT;
    end
  end

  assign when_PerformanceCounterPlugin_l271 = PerformanceCounterPlugin_logic_fsm_counterReaded[7];
  assign when_PerformanceCounterPlugin_l249 = (CsrAccessPlugin_bus_write_address[7] == 1'b0);
  assign when_PerformanceCounterPlugin_l255 = PerformanceCounterPlugin_logic_fsm_cmd_oh[1];
  assign PerformanceCounterPlugin_logic_fsm_onExit_BOOT = ((PerformanceCounterPlugin_logic_fsm_stateNext != PerformanceCounterPlugin_logic_fsm_BOOT) && (PerformanceCounterPlugin_logic_fsm_stateReg == PerformanceCounterPlugin_logic_fsm_BOOT));
  assign PerformanceCounterPlugin_logic_fsm_onExit_IDLE = ((PerformanceCounterPlugin_logic_fsm_stateNext != PerformanceCounterPlugin_logic_fsm_IDLE) && (PerformanceCounterPlugin_logic_fsm_stateReg == PerformanceCounterPlugin_logic_fsm_IDLE));
  assign PerformanceCounterPlugin_logic_fsm_onExit_READ_LOW = ((PerformanceCounterPlugin_logic_fsm_stateNext != PerformanceCounterPlugin_logic_fsm_READ_LOW) && (PerformanceCounterPlugin_logic_fsm_stateReg == PerformanceCounterPlugin_logic_fsm_READ_LOW));
  assign PerformanceCounterPlugin_logic_fsm_onExit_CALC_LOW = ((PerformanceCounterPlugin_logic_fsm_stateNext != PerformanceCounterPlugin_logic_fsm_CALC_LOW) && (PerformanceCounterPlugin_logic_fsm_stateReg == PerformanceCounterPlugin_logic_fsm_CALC_LOW));
  assign PerformanceCounterPlugin_logic_fsm_onExit_CSR_WRITE = ((PerformanceCounterPlugin_logic_fsm_stateNext != PerformanceCounterPlugin_logic_fsm_CSR_WRITE) && (PerformanceCounterPlugin_logic_fsm_stateReg == PerformanceCounterPlugin_logic_fsm_CSR_WRITE));
  assign PerformanceCounterPlugin_logic_fsm_onEntry_BOOT = ((PerformanceCounterPlugin_logic_fsm_stateNext == PerformanceCounterPlugin_logic_fsm_BOOT) && (PerformanceCounterPlugin_logic_fsm_stateReg != PerformanceCounterPlugin_logic_fsm_BOOT));
  assign PerformanceCounterPlugin_logic_fsm_onEntry_IDLE = ((PerformanceCounterPlugin_logic_fsm_stateNext == PerformanceCounterPlugin_logic_fsm_IDLE) && (PerformanceCounterPlugin_logic_fsm_stateReg != PerformanceCounterPlugin_logic_fsm_IDLE));
  assign PerformanceCounterPlugin_logic_fsm_onEntry_READ_LOW = ((PerformanceCounterPlugin_logic_fsm_stateNext == PerformanceCounterPlugin_logic_fsm_READ_LOW) && (PerformanceCounterPlugin_logic_fsm_stateReg != PerformanceCounterPlugin_logic_fsm_READ_LOW));
  assign PerformanceCounterPlugin_logic_fsm_onEntry_CALC_LOW = ((PerformanceCounterPlugin_logic_fsm_stateNext == PerformanceCounterPlugin_logic_fsm_CALC_LOW) && (PerformanceCounterPlugin_logic_fsm_stateReg != PerformanceCounterPlugin_logic_fsm_CALC_LOW));
  assign PerformanceCounterPlugin_logic_fsm_onEntry_CSR_WRITE = ((PerformanceCounterPlugin_logic_fsm_stateNext == PerformanceCounterPlugin_logic_fsm_CSR_WRITE) && (PerformanceCounterPlugin_logic_fsm_stateReg != PerformanceCounterPlugin_logic_fsm_CSR_WRITE));
  assign PerformanceCounterPlugin_logic_fsm_done = (PerformanceCounterPlugin_logic_fsm_stateReg == PerformanceCounterPlugin_logic_fsm_IDLE);
  always @(*) begin
    CsrAccessPlugin_logic_fsm_stateNext = CsrAccessPlugin_logic_fsm_stateReg;
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_READ : begin
        if(when_CsrAccessPlugin_l302) begin
          CsrAccessPlugin_logic_fsm_stateNext = CsrAccessPlugin_logic_fsm_WRITE;
        end
      end
      CsrAccessPlugin_logic_fsm_WRITE : begin
        if(when_CsrAccessPlugin_l331) begin
          CsrAccessPlugin_logic_fsm_stateNext = CsrAccessPlugin_logic_fsm_COMPLETION;
        end
      end
      CsrAccessPlugin_logic_fsm_COMPLETION : begin
        if(execute_ctrl2_down_isReady) begin
          CsrAccessPlugin_logic_fsm_stateNext = CsrAccessPlugin_logic_fsm_IDLE;
        end
      end
      default : begin
        if(CsrAccessPlugin_logic_fsm_inject_onDecodeDo) begin
          if(when_CsrAccessPlugin_l214) begin
            if(when_CsrAccessPlugin_l215) begin
              CsrAccessPlugin_logic_fsm_stateNext = CsrAccessPlugin_logic_fsm_READ;
            end
          end
          if(CsrAccessPlugin_logic_fsm_inject_sampled) begin
            if(!CsrAccessPlugin_logic_fsm_inject_trapReg) begin
              if(when_CsrAccessPlugin_l227) begin
                CsrAccessPlugin_logic_fsm_stateNext = CsrAccessPlugin_logic_fsm_READ;
              end
            end
          end
        end
      end
    endcase
    if(CsrAccessPlugin_logic_fsm_wantKill) begin
      CsrAccessPlugin_logic_fsm_stateNext = CsrAccessPlugin_logic_fsm_IDLE;
    end
  end

  assign when_CsrAccessPlugin_l302 = (! CsrAccessPlugin_bus_read_halt);
  assign when_CsrAccessPlugin_l331 = (! CsrAccessPlugin_bus_write_halt);
  assign when_CsrAccessPlugin_l214 = ((! CsrAccessPlugin_logic_fsm_inject_trap) && (! CsrAccessPlugin_bus_decode_trap));
  assign when_CsrAccessPlugin_l215 = (! CsrAccessPlugin_bus_decode_fence);
  assign when_CsrAccessPlugin_l227 = (! CsrAccessPlugin_bus_decode_fence);
  assign CsrAccessPlugin_logic_fsm_onExit_IDLE = ((CsrAccessPlugin_logic_fsm_stateNext != CsrAccessPlugin_logic_fsm_IDLE) && (CsrAccessPlugin_logic_fsm_stateReg == CsrAccessPlugin_logic_fsm_IDLE));
  assign CsrAccessPlugin_logic_fsm_onExit_READ = ((CsrAccessPlugin_logic_fsm_stateNext != CsrAccessPlugin_logic_fsm_READ) && (CsrAccessPlugin_logic_fsm_stateReg == CsrAccessPlugin_logic_fsm_READ));
  assign CsrAccessPlugin_logic_fsm_onExit_WRITE = ((CsrAccessPlugin_logic_fsm_stateNext != CsrAccessPlugin_logic_fsm_WRITE) && (CsrAccessPlugin_logic_fsm_stateReg == CsrAccessPlugin_logic_fsm_WRITE));
  assign CsrAccessPlugin_logic_fsm_onExit_COMPLETION = ((CsrAccessPlugin_logic_fsm_stateNext != CsrAccessPlugin_logic_fsm_COMPLETION) && (CsrAccessPlugin_logic_fsm_stateReg == CsrAccessPlugin_logic_fsm_COMPLETION));
  assign CsrAccessPlugin_logic_fsm_onEntry_IDLE = ((CsrAccessPlugin_logic_fsm_stateNext == CsrAccessPlugin_logic_fsm_IDLE) && (CsrAccessPlugin_logic_fsm_stateReg != CsrAccessPlugin_logic_fsm_IDLE));
  assign CsrAccessPlugin_logic_fsm_onEntry_READ = ((CsrAccessPlugin_logic_fsm_stateNext == CsrAccessPlugin_logic_fsm_READ) && (CsrAccessPlugin_logic_fsm_stateReg != CsrAccessPlugin_logic_fsm_READ));
  assign CsrAccessPlugin_logic_fsm_onEntry_WRITE = ((CsrAccessPlugin_logic_fsm_stateNext == CsrAccessPlugin_logic_fsm_WRITE) && (CsrAccessPlugin_logic_fsm_stateReg != CsrAccessPlugin_logic_fsm_WRITE));
  assign CsrAccessPlugin_logic_fsm_onEntry_COMPLETION = ((CsrAccessPlugin_logic_fsm_stateNext == CsrAccessPlugin_logic_fsm_COMPLETION) && (CsrAccessPlugin_logic_fsm_stateReg != CsrAccessPlugin_logic_fsm_COMPLETION));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      MmuPlugin_logic_satp_mode <= 4'b0000;
      MmuPlugin_logic_satp_ppn <= 44'h0;
      MmuPlugin_logic_status_mxr <= 1'b0;
      MmuPlugin_logic_status_sum <= 1'b0;
      PmpPlugin_logic_entries_0_address <= 21'h1fffff;
      PmpPlugin_logic_entries_0_cfg_read <= 1'b1;
      PmpPlugin_logic_entries_0_cfg_write <= 1'b1;
      PmpPlugin_logic_entries_0_cfg_execute <= 1'b1;
      PmpPlugin_logic_entries_0_cfg_kind <= 2'b11;
      PmpPlugin_logic_entries_0_cfg_locked <= 1'b0;
      PmpPlugin_logic_entries_1_address <= 21'h0;
      PmpPlugin_logic_entries_1_cfg_kind <= 2'b00;
      PmpPlugin_logic_entries_1_cfg_read <= 1'b0;
      PmpPlugin_logic_entries_1_cfg_write <= 1'b0;
      PmpPlugin_logic_entries_1_cfg_execute <= 1'b0;
      PmpPlugin_logic_entries_1_cfg_locked <= 1'b0;
      PmpPlugin_logic_entries_2_address <= 21'h0;
      PmpPlugin_logic_entries_2_cfg_kind <= 2'b00;
      PmpPlugin_logic_entries_2_cfg_read <= 1'b0;
      PmpPlugin_logic_entries_2_cfg_write <= 1'b0;
      PmpPlugin_logic_entries_2_cfg_execute <= 1'b0;
      PmpPlugin_logic_entries_2_cfg_locked <= 1'b0;
      PmpPlugin_logic_entries_3_address <= 21'h0;
      PmpPlugin_logic_entries_3_cfg_kind <= 2'b00;
      PmpPlugin_logic_entries_3_cfg_read <= 1'b0;
      PmpPlugin_logic_entries_3_cfg_write <= 1'b0;
      PmpPlugin_logic_entries_3_cfg_execute <= 1'b0;
      PmpPlugin_logic_entries_3_cfg_locked <= 1'b0;
      LsuL1Plugin_logic_refill_slots_0_valid <= 1'b0;
      LsuL1Plugin_logic_refill_slots_0_loaded <= 1'b1;
      LsuL1Plugin_logic_refill_pushCounter <= 32'h0;
      LsuL1Plugin_logic_refill_read_arbiter_lock <= 1'b0;
      LsuL1Plugin_logic_refill_read_wordIndex <= 3'b000;
      LsuL1Plugin_logic_refill_read_hadError <= 1'b0;
      LsuL1Plugin_logic_writeback_slots_0_valid <= 1'b0;
      LsuL1Plugin_logic_writeback_slots_0_busy <= 1'b0;
      LsuL1Plugin_logic_writeback_read_arbiter_lock <= 1'b0;
      LsuL1Plugin_logic_writeback_read_wordIndex <= 3'b000;
      LsuL1Plugin_logic_writeback_read_slotReadLast_valid <= 1'b0;
      LsuL1Plugin_logic_writeback_write_arbiter_lock <= 1'b0;
      LsuL1Plugin_logic_writeback_write_wordIndex <= 3'b000;
      LsuL1Plugin_logic_writeback_write_bufferRead_rValid <= 1'b0;
      LsuL1Plugin_logic_lsu_rb1_onBanks_0_busyReg <= 1'b0;
      LsuL1Plugin_logic_lsu_rb1_onBanks_1_busyReg <= 1'b0;
      LsuL1Plugin_logic_lsu_ctrl_hazardReg <= 1'b0;
      LsuL1Plugin_logic_lsu_ctrl_flushHazardReg <= 1'b0;
      LsuL1Plugin_logic_initializer_counter <= 7'h0;
      early0_MulPlugin_logic_writeback_buffer_valid <= 1'b0;
      early0_DivPlugin_logic_processing_cmdSent <= 1'b0;
      early0_DivPlugin_logic_processing_relaxer_hadRequest <= 1'b0;
      early0_DivPlugin_logic_processing_unscheduleRequest <= 1'b0;
      LsuL1Plugin_logic_bus_write_cmd_fork2_logic_linkEnable_0 <= 1'b1;
      LsuL1Plugin_logic_bus_write_cmd_fork2_logic_linkEnable_1 <= 1'b1;
      LsuL1Plugin_logic_bus_toAxi4_awRaw_payload_first <= 1'b1;
      LsuL1Plugin_logic_bus_toAxi4_awFiltred_rValid <= 1'b0;
      FetchL1Plugin_logic_invalidate_counter <= 7'h0;
      FetchL1Plugin_logic_invalidate_firstEver <= 1'b1;
      FetchL1Plugin_logic_refill_slots_0_valid <= 1'b0;
      FetchL1Plugin_logic_refill_slots_0_cmdSent <= 1'b1;
      FetchL1Plugin_logic_refill_pushCounter <= 32'h0;
      FetchL1Plugin_logic_refill_onCmd_locked <= 1'b0;
      FetchL1Plugin_logic_refill_onRsp_wordIndex <= 3'b000;
      FetchL1Plugin_logic_refill_onRsp_firstCycle <= 1'b1;
      FetchL1Plugin_logic_ctrl_plruLogic_buffer_regNext_valid <= 1'b0;
      FetchL1Plugin_logic_ctrl_trapSent <= 1'b0;
      FetchL1Plugin_logic_ctrl_firstCycle <= 1'b1;
      FetchL1Plugin_logic_ctrl_onEvents_waiting <= 1'b0;
      PrivilegedPlugin_logic_harts_0_privilege <= 2'b11;
      PrivilegedPlugin_logic_harts_0_m_status_mie <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_status_mpie <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_status_mpp <= 2'b00;
      PrivilegedPlugin_logic_harts_0_m_status_fs <= 2'b00;
      PrivilegedPlugin_logic_harts_0_m_status_tsr <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_status_tvm <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_status_tw <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_status_mprv <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_cause_interrupt <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_cause_code <= 4'b0000;
      PrivilegedPlugin_logic_harts_0_m_ip_meip <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_ip_mtip <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_ip_msip <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_ie_meie <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_ie_mtie <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_ie_msie <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_edeleg_iam <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_edeleg_bp <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_edeleg_eu <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_edeleg_es <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_edeleg_ipf <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_edeleg_lpf <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_edeleg_spf <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_ideleg_st <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_ideleg_se <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_ideleg_ss <= 1'b0;
      PrivilegedPlugin_logic_harts_0_s_cause_interrupt <= 1'b0;
      PrivilegedPlugin_logic_harts_0_s_cause_code <= 4'b0000;
      PrivilegedPlugin_logic_harts_0_s_status_sie <= 1'b0;
      PrivilegedPlugin_logic_harts_0_s_status_spie <= 1'b0;
      PrivilegedPlugin_logic_harts_0_s_status_spp <= 1'b0;
      PrivilegedPlugin_logic_harts_0_s_sstc_envcfg_enable <= 1'b0;
      PrivilegedPlugin_logic_harts_0_s_ip_seipSoft <= 1'b0;
      PrivilegedPlugin_logic_harts_0_s_ip_stipSoft <= 1'b0;
      PrivilegedPlugin_logic_harts_0_s_ip_ssip <= 1'b0;
      PrivilegedPlugin_logic_harts_0_s_ie_seie <= 1'b0;
      PrivilegedPlugin_logic_harts_0_s_ie_stie <= 1'b0;
      PrivilegedPlugin_logic_harts_0_s_ie_ssie <= 1'b0;
      BtbPlugin_logic_ras_ptr_push <= 2'b00;
      BtbPlugin_logic_ras_ptr_pop <= 2'b11;
      decode_ctrls_0_up_LANE_SEL_0_regNext <= 1'b0;
      PerformanceCounterPlugin_logic_ignoreNextCommit <= 1'b0;
      PerformanceCounterPlugin_logic_counters_cycle_value <= 8'h0;
      PerformanceCounterPlugin_logic_counters_cycle_mcounteren <= 1'b0;
      PerformanceCounterPlugin_logic_counters_cycle_scounteren <= 1'b0;
      PerformanceCounterPlugin_logic_counters_cycle_mcountinhibit <= 1'b0;
      PerformanceCounterPlugin_logic_counters_instret_value <= 8'h0;
      PerformanceCounterPlugin_logic_counters_instret_mcounteren <= 1'b0;
      PerformanceCounterPlugin_logic_counters_instret_scounteren <= 1'b0;
      PerformanceCounterPlugin_logic_counters_instret_mcountinhibit <= 1'b0;
      _zz_PerformanceCounterPlugin_logic_counters_instret_value <= 1'b0;
      LsuPlugin_logic_cbmCsr_menvcfg_cbie <= 2'b00;
      LsuPlugin_logic_cbmCsr_menvcfg_cbcfe <= 1'b0;
      LsuPlugin_logic_cbmCsr_senvcfg_cbie <= 2'b00;
      LsuPlugin_logic_cbmCsr_senvcfg_cbcfe <= 1'b0;
      LsuPlugin_logic_onAddress0_ls_storeId <= 12'h0;
      LsuPlugin_logic_onAddress0_access_waiter_valid <= 1'b0;
      execute_ctrl3_up_LsuL1_SEL_lane0 <= 1'b0;
      execute_ctrl4_up_LsuL1_SEL_lane0 <= 1'b0;
      LsuPlugin_logic_onCtrl_io_tooEarly <= 1'b0;
      LsuPlugin_logic_onCtrl_io_allowIt <= 1'b0;
      LsuPlugin_logic_onCtrl_io_doItReg <= 1'b0;
      LsuPlugin_logic_onCtrl_io_cmdSent <= 1'b0;
      LsuPlugin_logic_bus_rsp_toStream_rValid <= 1'b0;
      LsuPlugin_logic_onCtrl_rva_lrsc_reserved <= 1'b0;
      LsuPlugin_logic_onCtrl_fenceTrap_doItReg <= 1'b0;
      LsuPlugin_logic_onCtrl_cmbTrap_cmbTrigger <= 1'b0;
      LsuPlugin_logic_onCtrl_cmbTrap_pendingWritebacks <= 1'b0;
      LsuPlugin_logic_onCtrl_hartRegulation_valid <= 1'b0;
      LsuPlugin_logic_onCtrl_commitProbeToken <= 1'b0;
      AlignerPlugin_logic_feeder_harts_0_dopId <= 10'h0;
      AlignerPlugin_logic_buffer_mask <= 2'b00;
      AlignerPlugin_logic_buffer_last <= 2'b00;
      AlignerPlugin_logic_buffer_trap <= 1'b0;
      LsuCachelessAxi4Plugin_logic_bridge_tracker_pendings_0_valid <= 1'b0;
      LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_fork2_logic_linkEnable_0 <= 1'b1;
      LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_fork2_logic_linkEnable_1 <= 1'b1;
      DecoderPlugin_logic_harts_0_uopId <= 16'h0;
      DecoderPlugin_logic_interrupt_buffered <= 1'b0;
      decode_ctrls_1_up_LANE_SEL_0_regNext <= 1'b0;
      DispatchPlugin_logic_feeds_0_sent <= 1'b0;
      CsrRamPlugin_csrMapper_fired <= 1'b0;
      decode_ctrls_1_up_LANE_SEL_0_regNext_1 <= 1'b0;
      execute_ctrl0_down_LANE_SEL_lane0_regNext <= 1'b0;
      execute_ctrl2_down_LANE_SEL_lane0_regNext <= 1'b0;
      BtbPlugin_logic_applyIt_correctionSent <= 1'b0;
      decode_ctrls_1_up_LANE_SEL_0 <= 1'b0;
      TrapPlugin_logic_harts_0_interrupt_validBuffer <= 1'b0;
      TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidated <= 1'b0;
      TrapPlugin_logic_harts_0_trap_fsm_trapEnterDebug <= 1'b0;
      PcPlugin_logic_harts_0_self_id <= 10'h0;
      PcPlugin_logic_harts_0_self_increment <= 1'b0;
      PcPlugin_logic_harts_0_self_fault <= 1'b0;
      PcPlugin_logic_harts_0_self_state <= 39'h0000004000;
      PcPlugin_logic_harts_0_holdReg <= 1'b1;
      FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_value <= 1'b0;
      LsuPlugin_logic_translationStorage_logic_sl_0_allocId_value <= 2'b00;
      MmuPlugin_logic_refill_cacheRefillAny <= 1'b0;
      MmuPlugin_logic_accessBus_rsp_toStream_rValid <= 1'b0;
      MmuPlugin_logic_invalidate_busy <= 1'b0;
      HistoryPlugin_logic_onFetch_value <= 12'h0;
      PerformanceCounterPlugin_logic_interrupt_ip <= 1'b0;
      PerformanceCounterPlugin_logic_interrupt_ie <= 1'b0;
      PerformanceCounterPlugin_logic_interrupt_sup_deleg <= 1'b0;
      PerformanceCounterPlugin_logic_csrRead_fired <= 1'b0;
      PerformanceCounterPlugin_logic_csrWrite_fired <= 1'b0;
      CsrAccessPlugin_logic_fsm_inject_unfreeze <= 1'b0;
      CsrAccessPlugin_logic_fsm_inject_flushReg <= 1'b0;
      CsrAccessPlugin_logic_fsm_inject_sampled <= 1'b0;
      CsrRamPlugin_logic_readLogic_ohReg <= 3'b000;
      CsrRamPlugin_logic_readLogic_busy <= 1'b0;
      CsrRamPlugin_logic_flush_counter <= 5'h0;
      execute_ctrl1_up_LANE_SEL_lane0 <= 1'b0;
      execute_ctrl2_up_LANE_SEL_lane0 <= 1'b0;
      execute_ctrl3_up_LANE_SEL_lane0 <= 1'b0;
      execute_ctrl4_up_LANE_SEL_lane0 <= 1'b0;
      execute_ctrl5_up_LANE_SEL_lane0 <= 1'b0;
      integer_RegFilePlugin_logic_initalizer_counter <= 6'h0;
      _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_2 <= 60'h0;
      _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_2 <= 60'h0;
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_2 <= 60'h0;
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_2 <= 60'h0;
      _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_2 <= 60'h0;
      _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_2 <= 60'h0;
      fetch_logic_ctrls_1_up_valid <= 1'b0;
      fetch_logic_ctrls_2_up_valid <= 1'b0;
      decode_ctrls_1_up_valid <= 1'b0;
      LsuPlugin_logic_flusher_stateReg <= LsuPlugin_logic_flusher_IDLE;
      TrapPlugin_logic_harts_0_trap_fsm_stateReg <= TrapPlugin_logic_harts_0_trap_fsm_RESET;
      MmuPlugin_logic_refill_stateReg <= MmuPlugin_logic_refill_BOOT;
      PerformanceCounterPlugin_logic_fsm_stateReg <= PerformanceCounterPlugin_logic_fsm_BOOT;
      CsrAccessPlugin_logic_fsm_stateReg <= CsrAccessPlugin_logic_fsm_IDLE;
    end else begin
      if(when_PmpPlugin_l127) begin
        PmpPlugin_logic_entries_0_cfg_kind <= PmpPlugin_logic_entries_0_cfgNext_kind;
        PmpPlugin_logic_entries_0_cfg_read <= PmpPlugin_logic_entries_0_cfgNext_read;
        PmpPlugin_logic_entries_0_cfg_write <= PmpPlugin_logic_entries_0_cfgNext_write;
        PmpPlugin_logic_entries_0_cfg_execute <= PmpPlugin_logic_entries_0_cfgNext_execute;
        PmpPlugin_logic_entries_0_cfg_locked <= PmpPlugin_logic_entries_0_cfgNext_locked;
        if(when_PmpPlugin_l129) begin
          PmpPlugin_logic_entries_0_cfg_write <= 1'b0;
        end
      end
      if(when_PmpPlugin_l127_1) begin
        PmpPlugin_logic_entries_1_cfg_kind <= PmpPlugin_logic_entries_1_cfgNext_kind;
        PmpPlugin_logic_entries_1_cfg_read <= PmpPlugin_logic_entries_1_cfgNext_read;
        PmpPlugin_logic_entries_1_cfg_write <= PmpPlugin_logic_entries_1_cfgNext_write;
        PmpPlugin_logic_entries_1_cfg_execute <= PmpPlugin_logic_entries_1_cfgNext_execute;
        PmpPlugin_logic_entries_1_cfg_locked <= PmpPlugin_logic_entries_1_cfgNext_locked;
        if(when_PmpPlugin_l129_1) begin
          PmpPlugin_logic_entries_1_cfg_write <= 1'b0;
        end
      end
      if(when_PmpPlugin_l127_2) begin
        PmpPlugin_logic_entries_2_cfg_kind <= PmpPlugin_logic_entries_2_cfgNext_kind;
        PmpPlugin_logic_entries_2_cfg_read <= PmpPlugin_logic_entries_2_cfgNext_read;
        PmpPlugin_logic_entries_2_cfg_write <= PmpPlugin_logic_entries_2_cfgNext_write;
        PmpPlugin_logic_entries_2_cfg_execute <= PmpPlugin_logic_entries_2_cfgNext_execute;
        PmpPlugin_logic_entries_2_cfg_locked <= PmpPlugin_logic_entries_2_cfgNext_locked;
        if(when_PmpPlugin_l129_2) begin
          PmpPlugin_logic_entries_2_cfg_write <= 1'b0;
        end
      end
      if(when_PmpPlugin_l127_3) begin
        PmpPlugin_logic_entries_3_cfg_kind <= PmpPlugin_logic_entries_3_cfgNext_kind;
        PmpPlugin_logic_entries_3_cfg_read <= PmpPlugin_logic_entries_3_cfgNext_read;
        PmpPlugin_logic_entries_3_cfg_write <= PmpPlugin_logic_entries_3_cfgNext_write;
        PmpPlugin_logic_entries_3_cfg_execute <= PmpPlugin_logic_entries_3_cfgNext_execute;
        PmpPlugin_logic_entries_3_cfg_locked <= PmpPlugin_logic_entries_3_cfgNext_locked;
        if(when_PmpPlugin_l129_3) begin
          PmpPlugin_logic_entries_3_cfg_write <= 1'b0;
        end
      end
      if(LsuL1Plugin_logic_refill_slots_0_loadedSet) begin
        LsuL1Plugin_logic_refill_slots_0_loaded <= 1'b1;
      end
      if(LsuL1Plugin_logic_refill_slots_0_fire) begin
        LsuL1Plugin_logic_refill_slots_0_valid <= 1'b0;
      end
      if(LsuL1Plugin_logic_refill_push_valid) begin
        LsuL1Plugin_logic_refill_pushCounter <= (LsuL1Plugin_logic_refill_pushCounter + 32'h00000001);
      end
      if(when_LsuL1Plugin_l382) begin
        LsuL1Plugin_logic_refill_slots_0_valid <= 1'b1;
        LsuL1Plugin_logic_refill_slots_0_loaded <= 1'b0;
      end
      LsuL1Plugin_logic_refill_read_arbiter_lock <= LsuL1Plugin_logic_refill_read_arbiter_oh;
      if(LsuL1Plugin_logic_bus_read_cmd_fire) begin
        LsuL1Plugin_logic_refill_read_arbiter_lock <= 1'b0;
      end
      if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(LsuL1Plugin_logic_refill_read_writeReservation_win); // LsuL1Plugin.scala:L432
          `else
            if(!LsuL1Plugin_logic_refill_read_writeReservation_win) begin
              $display("FAILURE "); // LsuL1Plugin.scala:L432
              $finish;
            end
          `endif
        `endif
      end
      if(when_LsuL1Plugin_l453) begin
        LsuL1Plugin_logic_refill_read_hadError <= 1'b1;
      end
      if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(LsuL1Plugin_logic_refill_read_reservation_win); // LsuL1Plugin.scala:L462
          `else
            if(!LsuL1Plugin_logic_refill_read_reservation_win) begin
              $display("FAILURE "); // LsuL1Plugin.scala:L462
              $finish;
            end
          `endif
        `endif
        if(LsuL1Plugin_logic_refill_read_rspWithData) begin
          LsuL1Plugin_logic_refill_read_wordIndex <= (LsuL1Plugin_logic_refill_read_wordIndex + 3'b001);
        end
        if(when_LsuL1Plugin_l466) begin
          LsuL1Plugin_logic_refill_read_hadError <= 1'b0;
        end
      end
      if(LsuL1Plugin_logic_writeback_slots_0_fire) begin
        LsuL1Plugin_logic_writeback_slots_0_busy <= 1'b0;
      end
      if(when_LsuL1Plugin_l533) begin
        LsuL1Plugin_logic_writeback_slots_0_valid <= 1'b0;
      end
      if(when_LsuL1Plugin_l559) begin
        LsuL1Plugin_logic_writeback_slots_0_valid <= 1'b1;
        LsuL1Plugin_logic_writeback_slots_0_busy <= 1'b1;
      end
      LsuL1Plugin_logic_writeback_read_arbiter_lock <= LsuL1Plugin_logic_writeback_read_arbiter_oh;
      LsuL1Plugin_logic_writeback_read_wordIndex <= (LsuL1Plugin_logic_writeback_read_wordIndex + _zz_LsuL1Plugin_logic_writeback_read_wordIndex);
      if(when_LsuL1Plugin_l608) begin
        LsuL1Plugin_logic_writeback_read_arbiter_lock <= 1'b0;
      end
      LsuL1Plugin_logic_writeback_read_slotReadLast_valid <= LsuL1Plugin_logic_writeback_read_slotRead_valid;
      LsuL1Plugin_logic_writeback_write_arbiter_lock <= LsuL1Plugin_logic_writeback_write_arbiter_oh;
      LsuL1Plugin_logic_writeback_write_wordIndex <= (LsuL1Plugin_logic_writeback_write_wordIndex + _zz_LsuL1Plugin_logic_writeback_write_wordIndex);
      if(when_LsuL1Plugin_l679) begin
        LsuL1Plugin_logic_writeback_write_arbiter_lock <= 1'b0;
      end
      if(LsuL1Plugin_logic_writeback_write_bufferRead_ready) begin
        LsuL1Plugin_logic_writeback_write_bufferRead_rValid <= LsuL1Plugin_logic_writeback_write_bufferRead_valid;
      end
      if(LsuL1Plugin_logic_banks_0_usedByWriteback) begin
        LsuL1Plugin_logic_lsu_rb1_onBanks_0_busyReg <= 1'b1;
      end
      if(when_LsuL1Plugin_l738) begin
        LsuL1Plugin_logic_lsu_rb1_onBanks_0_busyReg <= 1'b0;
      end
      if(LsuL1Plugin_logic_banks_1_usedByWriteback) begin
        LsuL1Plugin_logic_lsu_rb1_onBanks_1_busyReg <= 1'b1;
      end
      if(when_LsuL1Plugin_l738_1) begin
        LsuL1Plugin_logic_lsu_rb1_onBanks_1_busyReg <= 1'b0;
      end
      LsuL1Plugin_logic_lsu_ctrl_hazardReg <= (execute_ctrl4_down_LsuL1_HAZARD_lane0 && execute_freeze_valid);
      LsuL1Plugin_logic_lsu_ctrl_flushHazardReg <= (execute_ctrl4_down_LsuL1_FLUSH_HAZARD_lane0 && execute_freeze_valid);
      if(execute_ctrl4_down_LsuL1_SEL_lane0) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert((_zz_56 <= 2'b01)); // LsuL1Plugin.scala:L904
          `else
            if(!(_zz_56 <= 2'b01)) begin
              $display("FAILURE Multiple way hit ???"); // LsuL1Plugin.scala:L904
              $finish;
            end
          `endif
        `endif
      end
      if(when_LsuL1Plugin_l926) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert((_zz_58 < 2'b10)); // LsuL1Plugin.scala:L927
          `else
            if(!(_zz_58 < 2'b10)) begin
              $display("FAILURE "); // LsuL1Plugin.scala:L927
              $finish;
            end
          `endif
        `endif
      end
      if(when_LsuL1Plugin_l1233) begin
        LsuL1Plugin_logic_initializer_counter <= (LsuL1Plugin_logic_initializer_counter + 7'h01);
      end
      early0_MulPlugin_logic_writeback_buffer_valid <= execute_freeze_valid;
      if(io_cmd_fire) begin
        early0_DivPlugin_logic_processing_cmdSent <= 1'b1;
      end
      if(execute_ctrl2_down_isReady) begin
        early0_DivPlugin_logic_processing_cmdSent <= 1'b0;
      end
      early0_DivPlugin_logic_processing_relaxer_hadRequest <= (early0_DivPlugin_logic_processing_request && execute_freeze_valid);
      early0_DivPlugin_logic_processing_unscheduleRequest <= execute_lane0_ctrls_2_upIsCancel;
      if(execute_ctrl2_down_isReady) begin
        early0_DivPlugin_logic_processing_unscheduleRequest <= 1'b0;
      end
      if(LsuL1Plugin_logic_bus_toAxi4_awRaw_fire) begin
        LsuL1Plugin_logic_bus_write_cmd_fork2_logic_linkEnable_0 <= 1'b0;
      end
      if(LsuL1Plugin_logic_bus_toAxi4_wRaw_fire) begin
        LsuL1Plugin_logic_bus_write_cmd_fork2_logic_linkEnable_1 <= 1'b0;
      end
      if(LsuL1Plugin_logic_bus_write_cmd_ready) begin
        LsuL1Plugin_logic_bus_write_cmd_fork2_logic_linkEnable_0 <= 1'b1;
        LsuL1Plugin_logic_bus_write_cmd_fork2_logic_linkEnable_1 <= 1'b1;
      end
      if(LsuL1Plugin_logic_bus_toAxi4_awRaw_fire) begin
        LsuL1Plugin_logic_bus_toAxi4_awRaw_payload_first <= LsuL1Plugin_logic_bus_toAxi4_awRaw_payload_last;
      end
      if(LsuL1Plugin_logic_bus_toAxi4_awFiltred_ready) begin
        LsuL1Plugin_logic_bus_toAxi4_awFiltred_rValid <= LsuL1Plugin_logic_bus_toAxi4_awFiltred_valid;
      end
      if(FetchL1Plugin_logic_invalidate_done) begin
        FetchL1Plugin_logic_invalidate_firstEver <= 1'b0;
      end
      if(when_FetchL1Plugin_l204) begin
        FetchL1Plugin_logic_invalidate_counter <= FetchL1Plugin_logic_invalidate_counterIncr;
      end
      if(when_FetchL1Plugin_l211) begin
        FetchL1Plugin_logic_invalidate_counter <= 7'h0;
      end
      if(when_FetchL1Plugin_l255) begin
        if(_zz_when_1) begin
          FetchL1Plugin_logic_refill_slots_0_valid <= 1'b1;
          FetchL1Plugin_logic_refill_slots_0_cmdSent <= 1'b0;
        end
        FetchL1Plugin_logic_refill_pushCounter <= (FetchL1Plugin_logic_refill_pushCounter + 32'h00000001);
      end
      if(FetchL1Plugin_logic_bus_cmd_valid) begin
        FetchL1Plugin_logic_refill_onCmd_locked <= 1'b1;
      end
      if(FetchL1Plugin_logic_bus_cmd_ready) begin
        FetchL1Plugin_logic_refill_onCmd_locked <= 1'b0;
      end
      if(FetchL1Plugin_logic_bus_cmd_ready) begin
        if(FetchL1Plugin_logic_refill_onCmd_oh[0]) begin
          FetchL1Plugin_logic_refill_slots_0_cmdSent <= 1'b1;
        end
      end
      if(FetchL1Plugin_logic_bus_rsp_fire) begin
        FetchL1Plugin_logic_refill_onRsp_firstCycle <= 1'b0;
      end
      if(FetchL1Plugin_logic_bus_rsp_valid) begin
        FetchL1Plugin_logic_refill_onRsp_wordIndex <= (FetchL1Plugin_logic_refill_onRsp_wordIndex + 3'b001);
        if(when_FetchL1Plugin_l330) begin
          FetchL1Plugin_logic_refill_onRsp_firstCycle <= 1'b1;
          FetchL1Plugin_logic_refill_slots_0_valid <= 1'b0;
        end
      end
      FetchL1Plugin_logic_ctrl_plruLogic_buffer_regNext_valid <= FetchL1Plugin_logic_ctrl_plruLogic_buffer_valid;
      if(FetchL1Plugin_logic_trapPort_valid) begin
        FetchL1Plugin_logic_ctrl_trapSent <= 1'b1;
      end
      if(fetch_logic_ctrls_2_up_isCancel) begin
        FetchL1Plugin_logic_ctrl_trapSent <= 1'b0;
      end
      if(fetch_logic_ctrls_2_up_isValid) begin
        FetchL1Plugin_logic_ctrl_firstCycle <= 1'b0;
      end
      if(when_FetchL1Plugin_l541) begin
        FetchL1Plugin_logic_ctrl_firstCycle <= 1'b1;
      end
      if(when_FetchL1Plugin_l549) begin
        FetchL1Plugin_logic_ctrl_onEvents_waiting <= 1'b0;
      end
      if(FetchL1Plugin_logic_events_miss) begin
        FetchL1Plugin_logic_ctrl_onEvents_waiting <= 1'b1;
      end
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert((! ((|FetchL1Plugin_logic_refill_slots_0_valid) && (! FetchL1Plugin_logic_invalidate_done)))); // FetchL1Plugin.scala:L556
        `else
          if(!(! ((|FetchL1Plugin_logic_refill_slots_0_valid) && (! FetchL1Plugin_logic_invalidate_done)))) begin
            $display("FAILURE "); // FetchL1Plugin.scala:L556
            $finish;
          end
        `endif
      `endif
      if(PrivilegedPlugin_logic_harts_0_xretAwayFromMachine) begin
        PrivilegedPlugin_logic_harts_0_m_status_mprv <= 1'b0;
      end
      PrivilegedPlugin_logic_harts_0_m_ip_meip <= PrivilegedPlugin_logic_harts_0_int_m_external;
      PrivilegedPlugin_logic_harts_0_m_ip_mtip <= PrivilegedPlugin_logic_harts_0_int_m_timer;
      PrivilegedPlugin_logic_harts_0_m_ip_msip <= PrivilegedPlugin_logic_harts_0_int_m_software;
      BtbPlugin_logic_ras_ptr_push <= (_zz_BtbPlugin_logic_ras_ptr_push - _zz_BtbPlugin_logic_ras_ptr_push_3);
      decode_ctrls_0_up_LANE_SEL_0_regNext <= decode_ctrls_0_up_LANE_SEL_0;
      if(when_CtrlLaneApi_l50) begin
        decode_ctrls_0_up_LANE_SEL_0_regNext <= 1'b0;
      end
      if(when_PerformanceCounterPlugin_l45) begin
        PerformanceCounterPlugin_logic_ignoreNextCommit <= 1'b0;
      end
      PerformanceCounterPlugin_logic_counters_cycle_value <= (PerformanceCounterPlugin_logic_counters_cycle_value + _zz_PerformanceCounterPlugin_logic_counters_cycle_value);
      _zz_PerformanceCounterPlugin_logic_counters_instret_value <= ((! PerformanceCounterPlugin_logic_counters_instret_mcountinhibit) ? PerformanceCounterPlugin_logic_commitCount : 1'b0);
      PerformanceCounterPlugin_logic_counters_instret_value <= (PerformanceCounterPlugin_logic_counters_instret_value + _zz_PerformanceCounterPlugin_logic_counters_instret_value_1);
      LsuPlugin_logic_onAddress0_ls_storeId <= (LsuPlugin_logic_onAddress0_ls_storeId + _zz_LsuPlugin_logic_onAddress0_ls_storeId);
      if(when_LsuPlugin_l264) begin
        LsuPlugin_logic_onAddress0_access_waiter_valid <= 1'b0;
      end
      LsuPlugin_logic_onCtrl_io_tooEarly <= 1'b1;
      if(execute_freeze_valid) begin
        LsuPlugin_logic_onCtrl_io_tooEarly <= 1'b0;
      end
      LsuPlugin_logic_onCtrl_io_allowIt <= 1'b0;
      if(when_LsuPlugin_l608) begin
        LsuPlugin_logic_onCtrl_io_allowIt <= 1'b1;
      end
      LsuPlugin_logic_onCtrl_io_doItReg <= LsuPlugin_logic_onCtrl_io_doIt;
      if(LsuPlugin_logic_bus_cmd_fire) begin
        LsuPlugin_logic_onCtrl_io_cmdSent <= 1'b1;
      end
      if(when_LsuPlugin_l612) begin
        LsuPlugin_logic_onCtrl_io_cmdSent <= 1'b0;
      end
      if(LsuPlugin_logic_bus_rsp_toStream_valid) begin
        LsuPlugin_logic_bus_rsp_toStream_rValid <= 1'b1;
      end
      if(LsuPlugin_logic_onCtrl_io_rsp_fire) begin
        LsuPlugin_logic_bus_rsp_toStream_rValid <= 1'b0;
      end
      if(when_LsuPlugin_l697) begin
        if(execute_ctrl4_down_LsuL1_STORE_lane0) begin
          LsuPlugin_logic_onCtrl_rva_lrsc_reserved <= 1'b0;
        end
      end
      if(when_LsuPlugin_l716) begin
        LsuPlugin_logic_onCtrl_rva_lrsc_reserved <= 1'b0;
      end
      if(when_LsuPlugin_l720) begin
        LsuPlugin_logic_onCtrl_rva_lrsc_reserved <= (! LsuPlugin_logic_onCtrl_rva_lrsc_reserved);
      end
      if(LsuPlugin_logic_onCtrl_fenceTrap_doIt) begin
        LsuPlugin_logic_onCtrl_fenceTrap_doItReg <= 1'b1;
      end
      if(when_LsuPlugin_l855) begin
        LsuPlugin_logic_onCtrl_fenceTrap_doItReg <= 1'b0;
      end
      if(when_LsuPlugin_l897) begin
        LsuPlugin_logic_onCtrl_cmbTrap_cmbTrigger <= ((execute_ctrl4_up_LANE_SEL_lane0 && execute_ctrl4_down_AguPlugin_SEL_lane0) && (execute_ctrl4_down_LsuL1_CLEAN_lane0 || execute_ctrl4_down_LsuL1_INVALID_lane0));
      end
      LsuPlugin_logic_onCtrl_cmbTrap_pendingWritebacks <= ((LsuPlugin_logic_onCtrl_cmbTrap_pendingWritebacks & (execute_freeze_valid ? 1'b1 : LsuL1_WRITEBACK_BUSY)) | (LsuPlugin_logic_onCtrl_cmbTrap_cmbTrigger ? LsuL1_WRITEBACK_BUSY : 1'b0));
      if(when_LsuPlugin_l986) begin
        if(when_LsuPlugin_l268) begin
          LsuPlugin_logic_onAddress0_access_waiter_valid <= 1'b1;
        end
      end
      if(when_LsuPlugin_l264_1) begin
        LsuPlugin_logic_onCtrl_hartRegulation_valid <= 1'b0;
      end
      if(when_LsuPlugin_l993) begin
        if(when_LsuPlugin_l268_1) begin
          LsuPlugin_logic_onCtrl_hartRegulation_valid <= 1'b1;
        end
      end
      if(LsuPlugin_logic_onCtrl_commitProbeReq) begin
        LsuPlugin_logic_onCtrl_commitProbeToken <= LsuPlugin_logic_onCtrl_lsuTrap;
      end
      if(when_AlignerPlugin_l171) begin
        AlignerPlugin_logic_feeder_harts_0_dopId <= (decode_ctrls_0_down_Decode_DOP_ID_0 + 10'h001);
      end
      if(AlignerPlugin_logic_buffer_downFire) begin
        AlignerPlugin_logic_buffer_mask <= (AlignerPlugin_logic_buffer_mask & (~ AlignerPlugin_logic_buffer_usedMask[1 : 0]));
        AlignerPlugin_logic_buffer_last <= (AlignerPlugin_logic_buffer_last & (~ AlignerPlugin_logic_buffer_usedMask[1 : 0]));
      end
      if(when_AlignerPlugin_l256) begin
        AlignerPlugin_logic_buffer_mask <= (fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK & (~ (AlignerPlugin_logic_buffer_downFire ? AlignerPlugin_logic_buffer_usedMask[3 : 2] : 2'b00)));
        AlignerPlugin_logic_buffer_trap <= fetch_logic_ctrls_2_down_TRAP;
        AlignerPlugin_logic_buffer_last <= fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_LAST;
      end
      if(LsuPlugin_logic_bus_rsp_valid) begin
        LsuCachelessAxi4Plugin_logic_bridge_tracker_pendings_0_valid <= 1'b0;
      end
      if(LsuPlugin_logic_bus_cmd_fire) begin
        LsuCachelessAxi4Plugin_logic_bridge_tracker_pendings_0_valid <= 1'b1;
      end
      if(LsuCachelessAxi4Plugin_logic_bridge_cmdFork_fire) begin
        LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_fork2_logic_linkEnable_0 <= 1'b0;
      end
      if(LsuCachelessAxi4Plugin_logic_bridge_dataFork_fire) begin
        LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_fork2_logic_linkEnable_1 <= 1'b0;
      end
      if(LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_ready) begin
        LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_fork2_logic_linkEnable_0 <= 1'b1;
        LsuCachelessAxi4Plugin_logic_bridge_cmdHalted_fork2_logic_linkEnable_1 <= 1'b1;
      end
      if(when_DecoderPlugin_l143) begin
        DecoderPlugin_logic_harts_0_uopId <= (DecoderPlugin_logic_harts_0_uopId + 16'h0001);
      end
      if(when_DecoderPlugin_l151) begin
        DecoderPlugin_logic_interrupt_buffered <= DecoderPlugin_logic_interrupt_async;
      end
      decode_ctrls_1_up_LANE_SEL_0_regNext <= decode_ctrls_1_up_LANE_SEL_0;
      if(when_CtrlLaneApi_l50_1) begin
        decode_ctrls_1_up_LANE_SEL_0_regNext <= 1'b0;
      end
      if(DispatchPlugin_logic_feeds_0_sending) begin
        DispatchPlugin_logic_feeds_0_sent <= 1'b1;
      end
      if(decode_ctrls_1_up_isMoving) begin
        DispatchPlugin_logic_feeds_0_sent <= 1'b0;
      end
      if(when_CsrRamPlugin_l97) begin
        CsrRamPlugin_csrMapper_fired <= 1'b1;
      end
      if(CsrAccessPlugin_bus_write_moving) begin
        CsrRamPlugin_csrMapper_fired <= 1'b0;
      end
      decode_ctrls_1_up_LANE_SEL_0_regNext_1 <= decode_ctrls_1_up_LANE_SEL_0;
      if(when_CtrlLaneApi_l50_2) begin
        decode_ctrls_1_up_LANE_SEL_0_regNext_1 <= 1'b0;
      end
      execute_ctrl0_down_LANE_SEL_lane0_regNext <= execute_ctrl0_down_LANE_SEL_lane0;
      if(when_CtrlLaneApi_l50_3) begin
        execute_ctrl0_down_LANE_SEL_lane0_regNext <= 1'b0;
      end
      execute_ctrl2_down_LANE_SEL_lane0_regNext <= execute_ctrl2_down_LANE_SEL_lane0;
      if(when_CtrlLaneApi_l50_4) begin
        execute_ctrl2_down_LANE_SEL_lane0_regNext <= 1'b0;
      end
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert((! (fetch_logic_ctrls_1_up_isValid && fetch_logic_ctrls_1_down_BtbPlugin_logic_readCmd_HAZARDS[0]))); // BtbPlugin.scala:L215
        `else
          if(!(! (fetch_logic_ctrls_1_up_isValid && fetch_logic_ctrls_1_down_BtbPlugin_logic_readCmd_HAZARDS[0]))) begin
            $display("FAILURE "); // BtbPlugin.scala:L215
            $finish;
          end
        `endif
      `endif
      if(fetch_logic_ctrls_1_up_isValid) begin
        BtbPlugin_logic_applyIt_correctionSent <= 1'b1;
      end
      if(when_BtbPlugin_l233) begin
        BtbPlugin_logic_applyIt_correctionSent <= 1'b0;
      end
      if(AlignerPlugin_logic_buffer_flushIt) begin
        AlignerPlugin_logic_buffer_mask <= 2'b00;
        AlignerPlugin_logic_buffer_last <= 2'b00;
      end
      TrapPlugin_logic_harts_0_interrupt_validBuffer <= TrapPlugin_logic_harts_0_interrupt_valid;
      if(TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidate_cmd_fire) begin
        TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidated <= 1'b1;
      end
      PcPlugin_logic_harts_0_holdReg <= PcPlugin_logic_harts_0_holdComb;
      PcPlugin_logic_harts_0_self_state <= PcPlugin_logic_harts_0_output_payload_pc;
      PcPlugin_logic_harts_0_self_fault <= PcPlugin_logic_harts_0_output_payload_fault;
      PcPlugin_logic_harts_0_self_increment <= 1'b0;
      if(PcPlugin_logic_harts_0_output_fire) begin
        PcPlugin_logic_harts_0_self_increment <= 1'b1;
        PcPlugin_logic_harts_0_self_state[1 : 1] <= 1'b0;
      end
      if(fetch_logic_ctrls_0_up_isFiring) begin
        PcPlugin_logic_harts_0_self_id <= (PcPlugin_logic_harts_0_self_id + 10'h001);
      end
      FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_value <= FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_valueNext;
      LsuPlugin_logic_translationStorage_logic_sl_0_allocId_value <= LsuPlugin_logic_translationStorage_logic_sl_0_allocId_valueNext;
      MmuPlugin_logic_refill_cacheRefillAny <= ((MmuPlugin_logic_refill_cacheRefillAny || MmuPlugin_logic_refill_cacheRefillAnySet) && (! 1'b0));
      if(MmuPlugin_logic_accessBus_rsp_toStream_ready) begin
        MmuPlugin_logic_accessBus_rsp_toStream_rValid <= MmuPlugin_logic_accessBus_rsp_toStream_valid;
      end
      if(when_MmuPlugin_l565) begin
        if(MmuPlugin_logic_invalidate_arbiter_io_output_valid) begin
          MmuPlugin_logic_invalidate_busy <= 1'b1;
        end
      end else begin
        if(when_MmuPlugin_l579) begin
          MmuPlugin_logic_invalidate_busy <= 1'b0;
        end
      end
      HistoryPlugin_logic_onFetch_value <= HistoryPlugin_logic_onFetch_valueNext;
      if(PerformanceCounterPlugin_logic_fsm_csrReadCmd_fire) begin
        PerformanceCounterPlugin_logic_csrRead_fired <= 1'b1;
      end
      if(CsrAccessPlugin_bus_read_moving) begin
        PerformanceCounterPlugin_logic_csrRead_fired <= 1'b0;
      end
      if(PerformanceCounterPlugin_logic_fsm_csrWriteCmd_fire) begin
        PerformanceCounterPlugin_logic_csrWrite_fired <= 1'b1;
      end
      if(CsrAccessPlugin_bus_write_moving) begin
        PerformanceCounterPlugin_logic_csrWrite_fired <= 1'b0;
      end
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert((! ((execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_down_CsrAccessPlugin_SEL_lane0) && execute_lane0_ctrls_2_upIsCancel))); // CsrAccessPlugin.scala:L137
        `else
          if(!(! ((execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_down_CsrAccessPlugin_SEL_lane0) && execute_lane0_ctrls_2_upIsCancel))) begin
            $display("FAILURE CsrAccessPlugin saw forbidden select && cancel request"); // CsrAccessPlugin.scala:L137
            $finish;
          end
        `endif
      `endif
      CsrAccessPlugin_logic_fsm_inject_unfreeze <= 1'b0;
      if(CsrAccessPlugin_logic_flushPort_valid) begin
        CsrAccessPlugin_logic_fsm_inject_flushReg <= 1'b1;
      end
      if(when_CsrAccessPlugin_l199) begin
        CsrAccessPlugin_logic_fsm_inject_flushReg <= 1'b0;
      end
      CsrAccessPlugin_logic_fsm_inject_sampled <= execute_freeze_valid;
      if(when_CsrAccessPlugin_l352) begin
        MmuPlugin_logic_status_mxr <= CsrAccessPlugin_bus_write_bits[19];
        MmuPlugin_logic_status_sum <= CsrAccessPlugin_bus_write_bits[18];
        PrivilegedPlugin_logic_harts_0_m_status_mpie <= CsrAccessPlugin_bus_write_bits[7];
        PrivilegedPlugin_logic_harts_0_m_status_mie <= CsrAccessPlugin_bus_write_bits[3];
        if(when_CsrService_l210) begin
          case(switch_PrivilegedPlugin_l581)
            2'b11 : begin
              PrivilegedPlugin_logic_harts_0_m_status_mpp <= 2'b11;
            end
            2'b01 : begin
              PrivilegedPlugin_logic_harts_0_m_status_mpp <= 2'b01;
            end
            2'b00 : begin
              PrivilegedPlugin_logic_harts_0_m_status_mpp <= 2'b00;
            end
            default : begin
            end
          endcase
        end
        PrivilegedPlugin_logic_harts_0_m_status_mprv <= CsrAccessPlugin_bus_write_bits[17];
        PrivilegedPlugin_logic_harts_0_m_status_fs <= CsrAccessPlugin_bus_write_bits[14 : 13];
        PrivilegedPlugin_logic_harts_0_m_status_tsr <= CsrAccessPlugin_bus_write_bits[22];
        PrivilegedPlugin_logic_harts_0_m_status_tvm <= CsrAccessPlugin_bus_write_bits[20];
        PrivilegedPlugin_logic_harts_0_m_status_tw <= CsrAccessPlugin_bus_write_bits[21];
        PrivilegedPlugin_logic_harts_0_s_status_spp <= CsrAccessPlugin_bus_write_bits[8 : 8];
        PrivilegedPlugin_logic_harts_0_s_status_spie <= CsrAccessPlugin_bus_write_bits[5];
        PrivilegedPlugin_logic_harts_0_s_status_sie <= CsrAccessPlugin_bus_write_bits[1];
      end
      if(when_CsrAccessPlugin_l352_1) begin
        MmuPlugin_logic_status_mxr <= CsrAccessPlugin_bus_write_bits[19];
        MmuPlugin_logic_status_sum <= CsrAccessPlugin_bus_write_bits[18];
        PrivilegedPlugin_logic_harts_0_s_status_spp <= CsrAccessPlugin_bus_write_bits[8 : 8];
        PrivilegedPlugin_logic_harts_0_s_status_spie <= CsrAccessPlugin_bus_write_bits[5];
        PrivilegedPlugin_logic_harts_0_s_status_sie <= CsrAccessPlugin_bus_write_bits[1];
        PrivilegedPlugin_logic_harts_0_m_status_fs <= CsrAccessPlugin_bus_write_bits[14 : 13];
      end
      if(when_CsrAccessPlugin_l359) begin
        if(when_CsrAccessPlugin_l352_2) begin
          MmuPlugin_logic_satp_mode <= CsrAccessPlugin_bus_write_bits[63 : 60];
          MmuPlugin_logic_satp_ppn <= CsrAccessPlugin_bus_write_bits[43 : 0];
        end
      end
      if(when_CsrAccessPlugin_l359_1) begin
        if(when_CsrAccessPlugin_l352_3) begin
          PmpPlugin_logic_entries_0_address[20 : 0] <= CsrAccessPlugin_bus_write_bits[29 : 9];
        end
      end
      if(when_CsrAccessPlugin_l359_2) begin
        if(when_CsrAccessPlugin_l352_5) begin
          PmpPlugin_logic_entries_1_address[20 : 0] <= CsrAccessPlugin_bus_write_bits[29 : 9];
        end
      end
      if(when_CsrAccessPlugin_l359_3) begin
        if(when_CsrAccessPlugin_l352_6) begin
          PmpPlugin_logic_entries_2_address[20 : 0] <= CsrAccessPlugin_bus_write_bits[29 : 9];
        end
      end
      if(when_CsrAccessPlugin_l359_4) begin
        if(when_CsrAccessPlugin_l352_7) begin
          PmpPlugin_logic_entries_3_address[20 : 0] <= CsrAccessPlugin_bus_write_bits[29 : 9];
        end
      end
      if(when_CsrAccessPlugin_l352_8) begin
        PrivilegedPlugin_logic_harts_0_m_cause_interrupt <= CsrAccessPlugin_bus_write_bits[63];
        PrivilegedPlugin_logic_harts_0_m_cause_code <= CsrAccessPlugin_bus_write_bits[3 : 0];
      end
      if(when_CsrAccessPlugin_l352_9) begin
        PrivilegedPlugin_logic_harts_0_s_ip_seipSoft <= CsrAccessPlugin_bus_write_bits[9];
        if(when_CsrService_l210) begin
          if(when_CsrService_l225) begin
            PrivilegedPlugin_logic_harts_0_s_ip_stipSoft <= CsrAccessPlugin_bus_write_bits[5];
          end
        end
        PrivilegedPlugin_logic_harts_0_s_ip_ssip <= CsrAccessPlugin_bus_write_bits[1];
        PerformanceCounterPlugin_logic_interrupt_ip <= CsrAccessPlugin_bus_write_bits[13];
      end
      if(when_CsrAccessPlugin_l352_10) begin
        PrivilegedPlugin_logic_harts_0_m_ie_meie <= CsrAccessPlugin_bus_write_bits[11];
        PrivilegedPlugin_logic_harts_0_m_ie_mtie <= CsrAccessPlugin_bus_write_bits[7];
        PrivilegedPlugin_logic_harts_0_m_ie_msie <= CsrAccessPlugin_bus_write_bits[3];
        PrivilegedPlugin_logic_harts_0_s_ie_seie <= CsrAccessPlugin_bus_write_bits[9];
        PrivilegedPlugin_logic_harts_0_s_ie_stie <= CsrAccessPlugin_bus_write_bits[5];
        PrivilegedPlugin_logic_harts_0_s_ie_ssie <= CsrAccessPlugin_bus_write_bits[1];
        PerformanceCounterPlugin_logic_interrupt_ie <= CsrAccessPlugin_bus_write_bits[13];
      end
      if(when_CsrAccessPlugin_l352_11) begin
        PrivilegedPlugin_logic_harts_0_m_edeleg_iam <= CsrAccessPlugin_bus_write_bits[0];
        PrivilegedPlugin_logic_harts_0_m_edeleg_bp <= CsrAccessPlugin_bus_write_bits[3];
        PrivilegedPlugin_logic_harts_0_m_edeleg_eu <= CsrAccessPlugin_bus_write_bits[8];
        PrivilegedPlugin_logic_harts_0_m_edeleg_es <= CsrAccessPlugin_bus_write_bits[9];
        PrivilegedPlugin_logic_harts_0_m_edeleg_ipf <= CsrAccessPlugin_bus_write_bits[12];
        PrivilegedPlugin_logic_harts_0_m_edeleg_lpf <= CsrAccessPlugin_bus_write_bits[13];
        PrivilegedPlugin_logic_harts_0_m_edeleg_spf <= CsrAccessPlugin_bus_write_bits[15];
      end
      if(when_CsrAccessPlugin_l352_12) begin
        PrivilegedPlugin_logic_harts_0_m_ideleg_se <= CsrAccessPlugin_bus_write_bits[9];
        PrivilegedPlugin_logic_harts_0_m_ideleg_st <= CsrAccessPlugin_bus_write_bits[5];
        PrivilegedPlugin_logic_harts_0_m_ideleg_ss <= CsrAccessPlugin_bus_write_bits[1];
        PerformanceCounterPlugin_logic_interrupt_sup_deleg <= CsrAccessPlugin_bus_write_bits[13];
      end
      if(when_CsrAccessPlugin_l352_13) begin
        PerformanceCounterPlugin_logic_counters_cycle_mcounteren <= CsrAccessPlugin_bus_write_bits[0];
        PerformanceCounterPlugin_logic_counters_instret_mcounteren <= CsrAccessPlugin_bus_write_bits[2];
      end
      if(when_CsrAccessPlugin_l352_14) begin
        PrivilegedPlugin_logic_harts_0_s_cause_interrupt <= CsrAccessPlugin_bus_write_bits[63];
        PrivilegedPlugin_logic_harts_0_s_cause_code <= CsrAccessPlugin_bus_write_bits[3 : 0];
      end
      if(when_CsrAccessPlugin_l352_15) begin
        if(when_CsrService_l210) begin
          if(PrivilegedPlugin_logic_harts_0_s_sstc_envcfg_allowUpdate) begin
            PrivilegedPlugin_logic_harts_0_s_sstc_envcfg_enable <= CsrAccessPlugin_bus_write_bits[63];
          end
        end
        LsuPlugin_logic_cbmCsr_menvcfg_cbie <= CsrAccessPlugin_bus_write_bits[5 : 4];
        LsuPlugin_logic_cbmCsr_menvcfg_cbcfe <= CsrAccessPlugin_bus_write_bits[6 : 6];
      end
      if(when_CsrAccessPlugin_l352_16) begin
        if(when_CsrService_l210) begin
          if(PrivilegedPlugin_logic_harts_0_m_ideleg_se) begin
            PrivilegedPlugin_logic_harts_0_s_ie_seie <= CsrAccessPlugin_bus_write_bits[9];
          end
        end
        if(when_CsrService_l210) begin
          if(PrivilegedPlugin_logic_harts_0_m_ideleg_st) begin
            PrivilegedPlugin_logic_harts_0_s_ie_stie <= CsrAccessPlugin_bus_write_bits[5];
          end
        end
        if(when_CsrService_l210) begin
          if(PrivilegedPlugin_logic_harts_0_m_ideleg_ss) begin
            PrivilegedPlugin_logic_harts_0_s_ie_ssie <= CsrAccessPlugin_bus_write_bits[1];
          end
        end
      end
      if(when_CsrAccessPlugin_l352_17) begin
        if(when_CsrService_l210) begin
          if(PrivilegedPlugin_logic_harts_0_m_ideleg_ss) begin
            PrivilegedPlugin_logic_harts_0_s_ip_ssip <= CsrAccessPlugin_bus_write_bits[1];
          end
        end
      end
      if(when_CsrAccessPlugin_l352_18) begin
        PerformanceCounterPlugin_logic_counters_cycle_scounteren <= CsrAccessPlugin_bus_write_bits[0];
        PerformanceCounterPlugin_logic_counters_instret_scounteren <= CsrAccessPlugin_bus_write_bits[2];
      end
      if(when_CsrAccessPlugin_l352_19) begin
        PerformanceCounterPlugin_logic_counters_cycle_mcountinhibit <= CsrAccessPlugin_bus_write_bits[0];
        PerformanceCounterPlugin_logic_counters_instret_mcountinhibit <= CsrAccessPlugin_bus_write_bits[2];
      end
      if(when_CsrAccessPlugin_l352_20) begin
        LsuPlugin_logic_cbmCsr_senvcfg_cbie <= CsrAccessPlugin_bus_write_bits[5 : 4];
        LsuPlugin_logic_cbmCsr_senvcfg_cbcfe <= CsrAccessPlugin_bus_write_bits[6 : 6];
      end
      CsrRamPlugin_logic_readLogic_ohReg <= (CsrRamPlugin_logic_readLogic_port_cmd_valid ? CsrRamPlugin_logic_readLogic_oh : 3'b000);
      CsrRamPlugin_logic_readLogic_busy <= CsrRamPlugin_logic_readLogic_port_cmd_valid;
      CsrRamPlugin_logic_flush_counter <= (CsrRamPlugin_logic_flush_counter + _zz_CsrRamPlugin_logic_flush_counter);
      if(when_RegFilePlugin_l132) begin
        integer_RegFilePlugin_logic_initalizer_counter <= (integer_RegFilePlugin_logic_initalizer_counter + 6'h01);
      end
      _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_2 <= _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_1;
      _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_2 <= _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_1;
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_2 <= _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_1;
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_2 <= _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_1;
      _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_2 <= _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_1;
      _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_2 <= _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_1;
      if(fetch_logic_ctrls_1_up_forgetOne) begin
        fetch_logic_ctrls_1_up_valid <= 1'b0;
      end
      if(fetch_logic_ctrls_0_down_isReady) begin
        fetch_logic_ctrls_1_up_valid <= fetch_logic_ctrls_0_down_isValid;
      end
      if(fetch_logic_ctrls_2_up_forgetOne) begin
        fetch_logic_ctrls_2_up_valid <= 1'b0;
      end
      if(fetch_logic_ctrls_1_down_isReady) begin
        fetch_logic_ctrls_2_up_valid <= fetch_logic_ctrls_1_down_isValid;
      end
      if(decode_ctrls_0_down_isReady) begin
        decode_ctrls_1_up_valid <= decode_ctrls_0_down_isValid;
      end
      if(decode_ctrls_0_down_isReady) begin
        decode_ctrls_1_up_LANE_SEL_0 <= decode_ctrls_0_down_LANE_SEL_0;
      end
      if(when_DecodePipelinePlugin_l70) begin
        decode_ctrls_1_up_LANE_SEL_0 <= 1'b0;
      end
      if(execute_ctrl0_down_isReady) begin
        execute_ctrl1_up_LANE_SEL_lane0 <= execute_ctrl0_down_LANE_SEL_lane0;
      end
      if(execute_ctrl1_down_isReady) begin
        execute_ctrl2_up_LANE_SEL_lane0 <= execute_ctrl1_down_LANE_SEL_lane0;
      end
      if(execute_ctrl2_down_isReady) begin
        execute_ctrl3_up_LANE_SEL_lane0 <= execute_ctrl2_down_LANE_SEL_lane0;
        execute_ctrl3_up_LsuL1_SEL_lane0 <= execute_ctrl2_down_LsuL1_SEL_lane0;
      end
      if(execute_ctrl3_down_isReady) begin
        execute_ctrl4_up_LANE_SEL_lane0 <= execute_ctrl3_down_LANE_SEL_lane0;
        execute_ctrl4_up_LsuL1_SEL_lane0 <= execute_ctrl3_down_LsuL1_SEL_lane0;
      end
      if(execute_ctrl4_down_isReady) begin
        execute_ctrl5_up_LANE_SEL_lane0 <= execute_ctrl4_down_LANE_SEL_lane0;
      end
      LsuPlugin_logic_flusher_stateReg <= LsuPlugin_logic_flusher_stateNext;
      TrapPlugin_logic_harts_0_trap_fsm_stateReg <= TrapPlugin_logic_harts_0_trap_fsm_stateNext;
      case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
        TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
        end
        TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
          TrapPlugin_logic_harts_0_trap_fsm_trapEnterDebug <= 1'b0;
          if(!when_TrapPlugin_l453) begin
            case(TrapPlugin_logic_harts_0_trap_pending_state_code)
              4'b0000 : begin
                `ifndef SYNTHESIS
                  `ifdef FORMAL
                    assert((! TrapPlugin_logic_harts_0_trap_fsm_buffer_i_valid)); // TrapPlugin.scala:L475
                  `else
                    if(!(! TrapPlugin_logic_harts_0_trap_fsm_buffer_i_valid)) begin
                      $display("FAILURE "); // TrapPlugin.scala:L475
                      $finish;
                    end
                  `endif
                `endif
              end
              4'b0001 : begin
              end
              4'b0010 : begin
              end
              4'b0100 : begin
              end
              4'b0101 : begin
              end
              4'b1000 : begin
              end
              4'b0110 : begin
              end
              4'b0111 : begin
              end
              default : begin
                `ifndef SYNTHESIS
                  `ifdef FORMAL
                    assert(1'b0); // TrapPlugin.scala:L528
                  `else
                    if(!1'b0) begin
                      $display("FAILURE Unexpected trap reason"); // TrapPlugin.scala:L528
                      $finish;
                    end
                  `endif
                `endif
              end
            endcase
          end
        end
        TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
        end
        TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
        end
        TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
        end
        TrapPlugin_logic_harts_0_trap_fsm_TRAP_WAIT : begin
        end
        TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
          PrivilegedPlugin_logic_harts_0_privilege <= TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_targetPrivilege;
          case(TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_targetPrivilege)
            2'b11 : begin
              PrivilegedPlugin_logic_harts_0_m_status_mie <= 1'b0;
              PrivilegedPlugin_logic_harts_0_m_status_mpie <= PrivilegedPlugin_logic_harts_0_m_status_mie;
              PrivilegedPlugin_logic_harts_0_m_status_mpp <= PrivilegedPlugin_logic_harts_0_privilege;
              PrivilegedPlugin_logic_harts_0_m_cause_code <= TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_code;
              PrivilegedPlugin_logic_harts_0_m_cause_interrupt <= TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_interrupt;
            end
            2'b01 : begin
              PrivilegedPlugin_logic_harts_0_s_status_sie <= 1'b0;
              PrivilegedPlugin_logic_harts_0_s_status_spie <= PrivilegedPlugin_logic_harts_0_s_status_sie;
              PrivilegedPlugin_logic_harts_0_s_status_spp <= PrivilegedPlugin_logic_harts_0_privilege[0 : 0];
              PrivilegedPlugin_logic_harts_0_s_cause_code <= TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_code;
              PrivilegedPlugin_logic_harts_0_s_cause_interrupt <= TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_interrupt;
            end
            default : begin
            end
          endcase
        end
        TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
        end
        TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
          PrivilegedPlugin_logic_harts_0_privilege <= TrapPlugin_logic_harts_0_trap_pending_xret_targetPrivilege;
          case(switch_TrapPlugin_l713)
            2'b11 : begin
              PrivilegedPlugin_logic_harts_0_m_status_mpp <= 2'b00;
              PrivilegedPlugin_logic_harts_0_m_status_mie <= PrivilegedPlugin_logic_harts_0_m_status_mpie;
              PrivilegedPlugin_logic_harts_0_m_status_mpie <= 1'b1;
            end
            2'b01 : begin
              PrivilegedPlugin_logic_harts_0_s_status_spp <= 1'b0;
              PrivilegedPlugin_logic_harts_0_s_status_sie <= PrivilegedPlugin_logic_harts_0_s_status_spie;
              PrivilegedPlugin_logic_harts_0_s_status_spie <= 1'b1;
            end
            default : begin
            end
          endcase
        end
        TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
        end
        TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
        end
        TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
        end
        TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
        end
        default : begin
        end
      endcase
      MmuPlugin_logic_refill_stateReg <= MmuPlugin_logic_refill_stateNext;
      PerformanceCounterPlugin_logic_fsm_stateReg <= PerformanceCounterPlugin_logic_fsm_stateNext;
      case(PerformanceCounterPlugin_logic_fsm_stateReg)
        PerformanceCounterPlugin_logic_fsm_IDLE : begin
        end
        PerformanceCounterPlugin_logic_fsm_READ_LOW : begin
        end
        PerformanceCounterPlugin_logic_fsm_CALC_LOW : begin
          if(when_PerformanceCounterPlugin_l271) begin
            if(_zz_PerformanceCounterPlugin_logic_fsm_cmd_address) begin
              PerformanceCounterPlugin_logic_counters_cycle_value[7] <= 1'b0;
            end
            if(_zz_PerformanceCounterPlugin_logic_fsm_cmd_address_1) begin
              PerformanceCounterPlugin_logic_counters_instret_value[7] <= 1'b0;
            end
          end
        end
        PerformanceCounterPlugin_logic_fsm_CSR_WRITE : begin
          if(when_PerformanceCounterPlugin_l249) begin
            if(_zz_PerformanceCounterPlugin_logic_fsm_cmd_address) begin
              PerformanceCounterPlugin_logic_counters_cycle_value <= _zz_PerformanceCounterPlugin_logic_counters_cycle_value_2[7:0];
              PerformanceCounterPlugin_logic_counters_cycle_value[7] <= 1'b0;
            end
            if(_zz_PerformanceCounterPlugin_logic_fsm_cmd_address_1) begin
              PerformanceCounterPlugin_logic_counters_instret_value <= _zz_PerformanceCounterPlugin_logic_counters_instret_value_2[7:0];
              PerformanceCounterPlugin_logic_counters_instret_value[7] <= 1'b0;
            end
          end
          if(when_PerformanceCounterPlugin_l255) begin
            PerformanceCounterPlugin_logic_ignoreNextCommit <= 1'b1;
          end
        end
        default : begin
        end
      endcase
      CsrAccessPlugin_logic_fsm_stateReg <= CsrAccessPlugin_logic_fsm_stateNext;
      case(CsrAccessPlugin_logic_fsm_stateReg)
        CsrAccessPlugin_logic_fsm_READ : begin
        end
        CsrAccessPlugin_logic_fsm_WRITE : begin
        end
        CsrAccessPlugin_logic_fsm_COMPLETION : begin
        end
        default : begin
          if(CsrAccessPlugin_logic_fsm_inject_onDecodeDo) begin
            if(CsrAccessPlugin_logic_fsm_inject_sampled) begin
              if(CsrAccessPlugin_logic_fsm_inject_trapReg) begin
                CsrAccessPlugin_logic_fsm_inject_unfreeze <= execute_freeze_valid;
              end
            end
          end
        end
      endcase
      case(CsrAccessPlugin_logic_fsm_stateNext)
        CsrAccessPlugin_logic_fsm_READ : begin
        end
        CsrAccessPlugin_logic_fsm_WRITE : begin
        end
        CsrAccessPlugin_logic_fsm_COMPLETION : begin
          CsrAccessPlugin_logic_fsm_inject_unfreeze <= 1'b1;
        end
        default : begin
        end
      endcase
      BtbPlugin_logic_ras_ptr_pop <= BtbPlugin_logic_ras_ptr_pop_aheadValue;
    end
  end

  always @(posedge clk) begin
    PmpPlugin_logic_entries_0_isNapot <= PmpPlugin_logic_entries_0_cfg_kind[1];
    PmpPlugin_logic_entries_0_isTor <= (PmpPlugin_logic_entries_0_cfg_kind == 2'b01);
    PmpPlugin_logic_entries_0_mask <= PmpPlugin_logic_entries_0_napot;
    PmpPlugin_logic_entries_1_isNapot <= PmpPlugin_logic_entries_1_cfg_kind[1];
    PmpPlugin_logic_entries_1_isTor <= (PmpPlugin_logic_entries_1_cfg_kind == 2'b01);
    PmpPlugin_logic_entries_1_mask <= PmpPlugin_logic_entries_1_napot;
    PmpPlugin_logic_entries_2_isNapot <= PmpPlugin_logic_entries_2_cfg_kind[1];
    PmpPlugin_logic_entries_2_isTor <= (PmpPlugin_logic_entries_2_cfg_kind == 2'b01);
    PmpPlugin_logic_entries_2_mask <= PmpPlugin_logic_entries_2_napot;
    PmpPlugin_logic_entries_3_isNapot <= PmpPlugin_logic_entries_3_cfg_kind[1];
    PmpPlugin_logic_entries_3_isTor <= (PmpPlugin_logic_entries_3_cfg_kind == 2'b01);
    PmpPlugin_logic_entries_3_mask <= PmpPlugin_logic_entries_3_napot;
    LsuL1Plugin_logic_refill_slots_0_loadedCounter <= (LsuL1Plugin_logic_refill_slots_0_loadedCounter + ((LsuL1Plugin_logic_refill_slots_0_loaded && (! LsuL1Plugin_logic_refill_slots_0_loadedDone)) && (! LsuL1Plugin_logic_slotsFreeze)));
    if(when_LsuL1Plugin_l386) begin
      LsuL1Plugin_logic_refill_slots_0_address <= LsuL1Plugin_logic_refill_push_payload_address;
      LsuL1Plugin_logic_refill_slots_0_way <= LsuL1Plugin_logic_refill_push_payload_way;
      LsuL1Plugin_logic_refill_slots_0_cmdSent <= 1'b0;
      LsuL1Plugin_logic_refill_slots_0_loadedCounter <= 1'b0;
      LsuL1Plugin_logic_refill_slots_0_victim <= LsuL1Plugin_logic_refill_push_payload_victim;
    end
    if(LsuL1Plugin_logic_refill_read_arbiter_oh[0]) begin
      if(LsuL1Plugin_logic_bus_read_cmd_ready) begin
        LsuL1Plugin_logic_refill_slots_0_cmdSent <= 1'b1;
      end
    end
    LsuL1Plugin_logic_writeback_slots_0_timer_counter <= (LsuL1Plugin_logic_writeback_slots_0_timer_counter + ((! LsuL1Plugin_logic_writeback_slots_0_timer_done) && (! LsuL1Plugin_logic_slotsFreeze)));
    if(when_LsuL1Plugin_l564) begin
      LsuL1Plugin_logic_writeback_slots_0_address <= LsuL1Plugin_logic_writeback_push_payload_address;
      LsuL1Plugin_logic_writeback_slots_0_way <= LsuL1Plugin_logic_writeback_push_payload_way;
      LsuL1Plugin_logic_writeback_slots_0_timer_counter <= 1'b0;
      LsuL1Plugin_logic_writeback_slots_0_writeCmdDone <= 1'b0;
      LsuL1Plugin_logic_writeback_slots_0_readCmdDone <= 1'b0;
      LsuL1Plugin_logic_writeback_slots_0_readRspDone <= 1'b0;
      LsuL1Plugin_logic_writeback_slots_0_victimBufferReady <= 1'b0;
    end
    if(when_LsuL1Plugin_l608) begin
      if(LsuL1Plugin_logic_writeback_read_arbiter_oh[0]) begin
        LsuL1Plugin_logic_writeback_slots_0_readCmdDone <= 1'b1;
      end
    end
    if(LsuL1Plugin_logic_writeback_read_slotRead_valid) begin
      LsuL1Plugin_logic_refill_slots_0_victim[0] <= 1'b0;
    end
    LsuL1Plugin_logic_writeback_read_slotReadLast_payload_last <= LsuL1Plugin_logic_writeback_read_slotRead_payload_last;
    LsuL1Plugin_logic_writeback_read_slotReadLast_payload_wordIndex <= LsuL1Plugin_logic_writeback_read_slotRead_payload_wordIndex;
    LsuL1Plugin_logic_writeback_read_slotReadLast_payload_way <= LsuL1Plugin_logic_writeback_read_slotRead_payload_way;
    if(LsuL1Plugin_logic_writeback_read_slotReadLast_valid) begin
      LsuL1Plugin_logic_writeback_slots_0_victimBufferReady <= 1'b1;
      if(LsuL1Plugin_logic_writeback_read_slotReadLast_payload_last) begin
        LsuL1Plugin_logic_writeback_slots_0_readRspDone <= 1'b1;
      end
    end
    if(when_LsuL1Plugin_l679) begin
      if(LsuL1Plugin_logic_writeback_write_arbiter_oh[0]) begin
        LsuL1Plugin_logic_writeback_slots_0_writeCmdDone <= 1'b1;
      end
    end
    if(LsuL1Plugin_logic_writeback_write_bufferRead_ready) begin
      LsuL1Plugin_logic_writeback_write_bufferRead_rData_address <= LsuL1Plugin_logic_writeback_write_bufferRead_payload_address;
      LsuL1Plugin_logic_writeback_write_bufferRead_rData_last <= LsuL1Plugin_logic_writeback_write_bufferRead_payload_last;
    end
    early0_MulPlugin_logic_writeback_buffer_data <= execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0[127 : 64];
    early0_DivPlugin_logic_processing_divRevertResult <= ((execute_ctrl2_down_RsUnsignedPlugin_RS1_REVERT_lane0 ^ (execute_ctrl2_down_RsUnsignedPlugin_RS2_REVERT_lane0 && (! execute_ctrl2_down_DivPlugin_REM_lane0))) && (! (((execute_ctrl2_down_RsUnsignedPlugin_RS2_FORMATED_lane0 == 64'h0) && execute_ctrl2_down_RsUnsignedPlugin_RS2_SIGNED_lane0) && (! execute_ctrl2_down_DivPlugin_REM_lane0))));
    early0_DivPlugin_logic_processing_a_delay_1 <= early0_DivPlugin_logic_processing_a;
    early0_DivPlugin_logic_processing_b_delay_1 <= early0_DivPlugin_logic_processing_b;
    if(LsuL1Plugin_logic_bus_toAxi4_awFiltred_ready) begin
      LsuL1Plugin_logic_bus_toAxi4_awFiltred_rData_last <= LsuL1Plugin_logic_bus_toAxi4_awFiltred_payload_last;
      LsuL1Plugin_logic_bus_toAxi4_awFiltred_rData_fragment_address <= LsuL1Plugin_logic_bus_toAxi4_awFiltred_payload_fragment_address;
      LsuL1Plugin_logic_bus_toAxi4_awFiltred_rData_fragment_data <= LsuL1Plugin_logic_bus_toAxi4_awFiltred_payload_fragment_data;
    end
    if(when_FetchL1Plugin_l255) begin
      if(_zz_when_1) begin
        FetchL1Plugin_logic_refill_slots_0_address <= FetchL1Plugin_logic_refill_start_address;
        FetchL1Plugin_logic_refill_slots_0_isIo <= FetchL1Plugin_logic_refill_start_isIo;
        FetchL1Plugin_logic_refill_slots_0_wayToAllocate <= FetchL1Plugin_logic_refill_start_wayToAllocate;
        FetchL1Plugin_logic_refill_slots_0_priority <= FetchL1Plugin_logic_refill_slots_0_valid;
      end
    end
    if(when_FetchL1Plugin_l276) begin
      FetchL1Plugin_logic_refill_onCmd_lockedOh <= FetchL1Plugin_logic_refill_onCmd_propoedOh;
    end
    FetchL1Plugin_logic_ctrl_plruLogic_buffer_regNext_payload_address <= FetchL1Plugin_logic_ctrl_plruLogic_buffer_payload_address;
    FetchL1Plugin_logic_ctrl_plruLogic_buffer_regNext_payload_data_0 <= FetchL1Plugin_logic_ctrl_plruLogic_buffer_payload_data_0;
    PrivilegedPlugin_logic_harts_0_s_ip_seipInput <= PrivilegedPlugin_logic_harts_0_int_s_external;
    if(BtbPlugin_logic_ras_readIt) begin
      BtbPlugin_logic_ras_read <= BtbPlugin_logic_ras_mem_stack_spinal_port0;
    end
    if(LsuPlugin_logic_onAddress0_flush_port_fire) begin
      LsuPlugin_logic_flusher_cmdCounter <= (LsuPlugin_logic_flusher_cmdCounter + 7'h01);
    end
    if(LsuPlugin_logic_bus_rsp_toStream_ready) begin
      LsuPlugin_logic_bus_rsp_toStream_rData_error <= LsuPlugin_logic_bus_rsp_toStream_payload_error;
      LsuPlugin_logic_bus_rsp_toStream_rData_data <= LsuPlugin_logic_bus_rsp_toStream_payload_data;
    end
    LsuPlugin_logic_onCtrl_rva_srcBuffer <= execute_ctrl4_down_LsuPlugin_logic_onCtrl_loadData_RESULT_lane0;
    LsuPlugin_logic_onCtrl_rva_aluBuffer <= LsuPlugin_logic_onCtrl_rva_alu_result;
    _zz_LsuPlugin_logic_onCtrl_rva_delay_0 <= (! execute_freeze_valid);
    _zz_LsuPlugin_logic_onCtrl_rva_delay_1 <= _zz_LsuPlugin_logic_onCtrl_rva_delay_0;
    if(when_LsuPlugin_l709) begin
      LsuPlugin_logic_onCtrl_rva_lrsc_age <= (LsuPlugin_logic_onCtrl_rva_lrsc_age + 6'h01);
    end
    if(when_LsuPlugin_l716) begin
      LsuPlugin_logic_onCtrl_rva_lrsc_age <= 6'h0;
    end
    if(when_LsuPlugin_l720) begin
      LsuPlugin_logic_onCtrl_rva_lrsc_address <= execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0;
      LsuPlugin_logic_onCtrl_rva_lrsc_age <= 6'h0;
    end
    if(when_LsuPlugin_l949) begin
      LsuPlugin_logic_flusher_cmdCounter <= {1'd0, _zz_LsuPlugin_logic_flusher_cmdCounter};
    end
    if(when_LsuPlugin_l986) begin
      if(when_LsuPlugin_l268) begin
        LsuPlugin_logic_onAddress0_access_waiter_refill <= execute_ctrl4_down_LsuL1_WAIT_REFILL_lane0;
      end
    end
    if(when_LsuPlugin_l993) begin
      if(when_LsuPlugin_l268_1) begin
        LsuPlugin_logic_onCtrl_hartRegulation_refill <= execute_ctrl4_down_LsuL1_WAIT_REFILL_lane0;
      end
    end
    if(when_AlignerPlugin_l256) begin
      AlignerPlugin_logic_buffer_data <= fetch_logic_ctrls_2_down_Fetch_WORD;
      AlignerPlugin_logic_buffer_pc <= fetch_logic_ctrls_2_down_Fetch_WORD_PC;
      AlignerPlugin_logic_buffer_hm_Fetch_ID <= fetch_logic_ctrls_2_down_Fetch_ID;
      AlignerPlugin_logic_buffer_hm_GSharePlugin_GSHARE_COUNTER_0 <= fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_0;
      AlignerPlugin_logic_buffer_hm_GSharePlugin_GSHARE_COUNTER_1 <= fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_1;
      AlignerPlugin_logic_buffer_hm_Prediction_BRANCH_HISTORY <= fetch_logic_ctrls_2_down_Prediction_BRANCH_HISTORY;
      AlignerPlugin_logic_buffer_hm_Prediction_WORD_SLICES_BRANCH <= fetch_logic_ctrls_2_down_Prediction_WORD_SLICES_BRANCH;
      AlignerPlugin_logic_buffer_hm_Prediction_WORD_SLICES_TAKEN <= fetch_logic_ctrls_2_down_Prediction_WORD_SLICES_TAKEN;
      AlignerPlugin_logic_buffer_hm_Prediction_WORD_JUMP_PC <= fetch_logic_ctrls_2_down_Prediction_WORD_JUMP_PC;
      AlignerPlugin_logic_buffer_hm_Prediction_WORD_JUMPED <= fetch_logic_ctrls_2_down_Prediction_WORD_JUMPED;
      AlignerPlugin_logic_buffer_hm_Prediction_WORD_JUMP_SLICE <= fetch_logic_ctrls_2_down_Prediction_WORD_JUMP_SLICE;
    end
    if(LsuPlugin_logic_bus_cmd_fire) begin
      LsuCachelessAxi4Plugin_logic_bridge_tracker_pendings_0_hash <= LsuCachelessAxi4Plugin_logic_bridge_cmdHash;
      LsuCachelessAxi4Plugin_logic_bridge_tracker_pendings_0_mask <= LsuPlugin_logic_bus_cmd_payload_mask;
      LsuCachelessAxi4Plugin_logic_bridge_tracker_pendings_0_io <= LsuPlugin_logic_bus_cmd_payload_io;
    end
    TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_triggered_id <= (_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_triggered_id_1 ? (_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_triggered_id ? TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_0_id : TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_1_id) : TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_2_id);
    TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_triggered_priority <= (_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_triggered_id_1 ? _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_triggered_priority : TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_2_priority);
    TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_triggered_privilege <= (_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_triggered_id_1 ? _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_triggered_privilege : TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_2_privilege);
    TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_triggered_valid <= (_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_triggered_id_1 ? _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_triggered_valid : TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_0_interrupts_2_valid);
    TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id <= (_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_10 ? (_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_9 ? (_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id ? TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_0_id : TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_1_id) : (_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_4 ? TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_2_id : TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_3_id)) : (_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_8 ? TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_4_id : TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_interrupts_5_id));
    TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_priority <= (_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_10 ? _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_priority_1 : _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_priority);
    TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_privilege <= (_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_10 ? _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_privilege_1 : _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_privilege);
    TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_valid <= (_zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_id_10 ? _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_valid_1 : _zz_TrapPlugin_logic_harts_0_interrupt_privilegeTriggers_1_triggered_valid);
    if(TrapPlugin_logic_harts_0_trap_pending_arbiter_down_valid) begin
      TrapPlugin_logic_harts_0_trap_pending_state_exception <= TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception;
      TrapPlugin_logic_harts_0_trap_pending_state_tval <= TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_tval;
      TrapPlugin_logic_harts_0_trap_pending_state_code <= TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_code;
      TrapPlugin_logic_harts_0_trap_pending_state_arg <= TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_arg;
    end
    if(TrapPlugin_logic_harts_0_trap_trigger_valid) begin
      TrapPlugin_logic_harts_0_trap_pending_pc <= execute_ctrl4_down_PC_lane0;
      TrapPlugin_logic_harts_0_trap_pending_history <= execute_ctrl4_down_Prediction_BRANCH_HISTORY_lane0;
      TrapPlugin_logic_harts_0_trap_pending_slices <= (_zz_TrapPlugin_logic_harts_0_trap_pending_slices + 2'b01);
    end
    if(TrapPlugin_logic_harts_0_trap_fsm_buffer_sampleIt) begin
      TrapPlugin_logic_harts_0_trap_fsm_buffer_i_valid <= TrapPlugin_logic_harts_0_interrupt_valid;
    end
    if(TrapPlugin_logic_harts_0_trap_fsm_buffer_sampleIt) begin
      TrapPlugin_logic_harts_0_trap_fsm_buffer_i_code <= TrapPlugin_logic_harts_0_interrupt_code;
    end
    if(TrapPlugin_logic_harts_0_trap_fsm_buffer_sampleIt) begin
      TrapPlugin_logic_harts_0_trap_fsm_buffer_i_targetPrivilege <= TrapPlugin_logic_harts_0_interrupt_targetPrivilege;
    end
    TrapPlugin_logic_harts_0_trap_fsm_jumpTarget <= (TrapPlugin_logic_harts_0_trap_pending_pc + _zz_TrapPlugin_logic_harts_0_trap_fsm_jumpTarget);
    if(when_TrapPlugin_l602) begin
      TrapPlugin_logic_harts_0_trap_fsm_readed <= TrapPlugin_logic_harts_0_crsPorts_read_data;
    end
    if(MmuPlugin_logic_accessBus_rsp_toStream_ready) begin
      MmuPlugin_logic_accessBus_rsp_toStream_rData_data <= MmuPlugin_logic_accessBus_rsp_toStream_payload_data;
      MmuPlugin_logic_accessBus_rsp_toStream_rData_error <= MmuPlugin_logic_accessBus_rsp_toStream_payload_error;
      MmuPlugin_logic_accessBus_rsp_toStream_rData_redo <= MmuPlugin_logic_accessBus_rsp_toStream_payload_redo;
      MmuPlugin_logic_accessBus_rsp_toStream_rData_waitAny <= MmuPlugin_logic_accessBus_rsp_toStream_payload_waitAny;
    end
    if(when_MmuPlugin_l565) begin
      MmuPlugin_logic_invalidate_counter <= 5'h0;
    end else begin
      MmuPlugin_logic_invalidate_counter <= (MmuPlugin_logic_invalidate_counter + 5'h01);
    end
    _zz_PerformanceCounterPlugin_logic_events_sums_0 <= early0_BranchPlugin_logic_events_branchMiss;
    _zz_PerformanceCounterPlugin_logic_events_sums_1 <= early0_BranchPlugin_logic_events_branchCount;
    _zz_PerformanceCounterPlugin_logic_events_sums_2 <= LsuPlugin_logic_events_waiting;
    _zz_PerformanceCounterPlugin_logic_events_sums_3 <= LsuL1Plugin_logic_events_loadAccess;
    _zz_PerformanceCounterPlugin_logic_events_sums_4 <= LsuL1Plugin_logic_events_loadMiss;
    _zz_PerformanceCounterPlugin_logic_events_sums_5 <= FetchL1Plugin_logic_events_access;
    _zz_PerformanceCounterPlugin_logic_events_sums_6 <= FetchL1Plugin_logic_events_miss;
    _zz_PerformanceCounterPlugin_logic_events_sums_7 <= FetchL1Plugin_logic_events_waiting;
    _zz_PerformanceCounterPlugin_logic_events_sums_8 <= PerformanceCounterPlugin_logic_eventCycles;
    _zz_PerformanceCounterPlugin_logic_events_sums_9 <= PerformanceCounterPlugin_logic_eventInstructions_0;
    _zz_PerformanceCounterPlugin_logic_events_sums_10 <= DispatchPlugin_logic_events_frontendStall;
    _zz_PerformanceCounterPlugin_logic_events_sums_11 <= DispatchPlugin_logic_events_backendStall;
    _zz_PerformanceCounterPlugin_logic_events_sums_12 <= MmuPlugin_logic_refill_events_onStorage_0_waiting;
    _zz_PerformanceCounterPlugin_logic_events_sums_13 <= MmuPlugin_logic_refill_events_onStorage_1_waiting;
    CsrAccessPlugin_logic_fsm_interface_read <= ((execute_ctrl2_down_CsrAccessPlugin_SEL_lane0 && (! CsrAccessPlugin_logic_fsm_inject_trap)) && CsrAccessPlugin_logic_fsm_inject_csrRead);
    CsrAccessPlugin_logic_fsm_interface_write <= ((execute_ctrl2_down_CsrAccessPlugin_SEL_lane0 && (! CsrAccessPlugin_logic_fsm_inject_trap)) && CsrAccessPlugin_logic_fsm_inject_csrWrite);
    CsrAccessPlugin_logic_fsm_inject_trapReg <= CsrAccessPlugin_logic_fsm_inject_trap;
    CsrAccessPlugin_logic_fsm_inject_busTrapReg <= CsrAccessPlugin_bus_decode_trap;
    CsrAccessPlugin_logic_fsm_inject_busTrapCodeReg <= CsrAccessPlugin_bus_decode_trapCode;
    CsrAccessPlugin_logic_fsm_interface_onWriteBits <= CsrAccessPlugin_logic_fsm_writeLogic_alu_result;
    if(when_CsrAccessPlugin_l352_13) begin
      PrivilegedPlugin_logic_harts_0_mcounteren_tm <= CsrAccessPlugin_bus_write_bits[1];
    end
    if(fetch_logic_ctrls_0_down_isReady) begin
      fetch_logic_ctrls_1_up_Fetch_WORD_PC <= fetch_logic_ctrls_0_down_Fetch_WORD_PC;
      fetch_logic_ctrls_1_up_Fetch_PC_FAULT <= fetch_logic_ctrls_0_down_Fetch_PC_FAULT;
      fetch_logic_ctrls_1_up_Fetch_ID <= fetch_logic_ctrls_0_down_Fetch_ID;
      _zz_1 <= 1'b0;
      fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_PLRU_BYPASS_VALID <= fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_VALID;
      fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_0 <= fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_0;
      fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_TAGS_UPDATE <= fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE;
      fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_TAGS_UPDATE_ADDRESS <= fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE_ADDRESS;
      fetch_logic_ctrls_1_up_GSharePlugin_logic_HASH <= fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH;
      fetch_logic_ctrls_1_up_Prediction_BRANCH_HISTORY <= fetch_logic_ctrls_0_down_Prediction_BRANCH_HISTORY;
      fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_valid <= fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_valid;
      fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_address <= fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_address;
      fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_data_0 <= fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_data_0;
      fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_data_1 <= fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_data_1;
      fetch_logic_ctrls_1_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_PERM_OK <= fetch_logic_ctrls_0_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_PERM_OK;
      fetch_logic_ctrls_1_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_PERM_OK <= fetch_logic_ctrls_0_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_PERM_OK;
      fetch_logic_ctrls_1_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_PERM_OK <= fetch_logic_ctrls_0_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_PERM_OK;
      fetch_logic_ctrls_1_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_PERM_OK <= fetch_logic_ctrls_0_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_PERM_OK;
      fetch_logic_ctrls_1_up_FetchL1Plugin_logic_pmpPort_logic_NEED_HIT <= fetch_logic_ctrls_0_down_FetchL1Plugin_logic_pmpPort_logic_NEED_HIT;
      fetch_logic_ctrls_1_up_BtbPlugin_logic_readCmd_HAZARDS <= fetch_logic_ctrls_0_down_BtbPlugin_logic_readCmd_HAZARDS;
    end
    if(fetch_logic_ctrls_1_down_isReady) begin
      fetch_logic_ctrls_2_up_Fetch_WORD_PC <= fetch_logic_ctrls_1_down_Fetch_WORD_PC;
      fetch_logic_ctrls_2_up_Fetch_PC_FAULT <= fetch_logic_ctrls_1_down_Fetch_PC_FAULT;
      fetch_logic_ctrls_2_up_Fetch_ID <= fetch_logic_ctrls_1_down_Fetch_ID;
      fetch_logic_ctrls_2_up_Prediction_BRANCH_HISTORY <= fetch_logic_ctrls_1_down_Prediction_BRANCH_HISTORY;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_PERM_OK <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_PERM_OK;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_PERM_OK <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_PERM_OK;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_PERM_OK <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_PERM_OK;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_PERM_OK <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_PERM_OK;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_pmpPort_logic_NEED_HIT <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_NEED_HIT;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_0_loaded <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_loaded;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_0_error <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_error;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_0_address <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_address;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_1_loaded <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_loaded;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_1_error <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_error;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_1_address <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_address;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_PLRU_BYPASSED_0 <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_PLRU_BYPASSED_0;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_BANKS_MUXES_0 <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_0;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_BANKS_MUXES_1 <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_1;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_HAZARD <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_HAZARD;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_HITS_0 <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HITS_0;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_HITS_1 <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HITS_1;
      fetch_logic_ctrls_2_up_MMU_BYPASS_TRANSLATION <= fetch_logic_ctrls_1_down_MMU_BYPASS_TRANSLATION;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_HIT <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HIT;
      fetch_logic_ctrls_2_up_GSharePlugin_GSHARE_COUNTER_0 <= fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0;
      fetch_logic_ctrls_2_up_GSharePlugin_GSHARE_COUNTER_1 <= fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_1;
      fetch_logic_ctrls_2_up_MMU_TRANSLATED <= fetch_logic_ctrls_1_down_MMU_TRANSLATED;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_napot_HIT <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_napot_HIT;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_tor_BIGGER <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_0_tor_BIGGER;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_napot_HIT <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_napot_HIT;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_tor_BIGGER <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_1_tor_BIGGER;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_napot_HIT <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_napot_HIT;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_tor_BIGGER <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_2_tor_BIGGER;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_napot_HIT <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_napot_HIT;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_tor_BIGGER <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_pmpPort_logic_onEntries_3_tor_BIGGER;
      fetch_logic_ctrls_2_up_Prediction_WORD_JUMPED <= fetch_logic_ctrls_1_down_Prediction_WORD_JUMPED;
      fetch_logic_ctrls_2_up_Prediction_WORD_JUMP_SLICE <= fetch_logic_ctrls_1_down_Prediction_WORD_JUMP_SLICE;
      fetch_logic_ctrls_2_up_Prediction_WORD_JUMP_PC <= fetch_logic_ctrls_1_down_Prediction_WORD_JUMP_PC;
      fetch_logic_ctrls_2_up_Prediction_WORD_SLICES_BRANCH <= fetch_logic_ctrls_1_down_Prediction_WORD_SLICES_BRANCH;
      fetch_logic_ctrls_2_up_Prediction_WORD_SLICES_TAKEN <= fetch_logic_ctrls_1_down_Prediction_WORD_SLICES_TAKEN;
      fetch_logic_ctrls_2_up_MMU_HAZARD <= fetch_logic_ctrls_1_down_MMU_HAZARD;
      fetch_logic_ctrls_2_up_MMU_REFILL <= fetch_logic_ctrls_1_down_MMU_REFILL;
      fetch_logic_ctrls_2_up_MMU_ALLOW_EXECUTE <= fetch_logic_ctrls_1_down_MMU_ALLOW_EXECUTE;
      fetch_logic_ctrls_2_up_MMU_PAGE_FAULT <= fetch_logic_ctrls_1_down_MMU_PAGE_FAULT;
      fetch_logic_ctrls_2_up_MMU_ACCESS_FAULT <= fetch_logic_ctrls_1_down_MMU_ACCESS_FAULT;
    end
    if(decode_ctrls_0_down_isReady) begin
      decode_ctrls_1_up_Decode_INSTRUCTION_0 <= decode_ctrls_0_down_Decode_INSTRUCTION_0;
      decode_ctrls_1_up_Decode_DECOMPRESSION_FAULT_0 <= decode_ctrls_0_down_Decode_DECOMPRESSION_FAULT_0;
      decode_ctrls_1_up_Decode_INSTRUCTION_RAW_0 <= decode_ctrls_0_down_Decode_INSTRUCTION_RAW_0;
      decode_ctrls_1_up_Decode_INSTRUCTION_SLICE_COUNT_0 <= decode_ctrls_0_down_Decode_INSTRUCTION_SLICE_COUNT_0;
      decode_ctrls_1_up_PC_0 <= decode_ctrls_0_down_PC_0;
      decode_ctrls_1_up_Decode_DOP_ID_0 <= decode_ctrls_0_down_Decode_DOP_ID_0;
      decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_0_0 <= decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_0_0;
      decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_0_1 <= decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_0_1;
      decode_ctrls_1_up_Prediction_BRANCH_HISTORY_0 <= decode_ctrls_0_down_Prediction_BRANCH_HISTORY_0;
      decode_ctrls_1_up_TRAP_0 <= decode_ctrls_0_down_TRAP_0;
      decode_ctrls_1_up_Prediction_ALIGNED_JUMPED_0 <= decode_ctrls_0_down_Prediction_ALIGNED_JUMPED_0;
      decode_ctrls_1_up_Prediction_ALIGNED_JUMPED_PC_0 <= decode_ctrls_0_down_Prediction_ALIGNED_JUMPED_PC_0;
      decode_ctrls_1_up_Prediction_ALIGNED_SLICES_BRANCH_0 <= decode_ctrls_0_down_Prediction_ALIGNED_SLICES_BRANCH_0;
      decode_ctrls_1_up_Prediction_ALIGNED_SLICES_TAKEN_0 <= decode_ctrls_0_down_Prediction_ALIGNED_SLICES_TAKEN_0;
      decode_ctrls_1_up_Prediction_ALIGN_REDO_0 <= decode_ctrls_0_down_Prediction_ALIGN_REDO_0;
    end
    if(execute_ctrl0_down_isReady) begin
      execute_ctrl1_up_Decode_UOP_lane0 <= execute_ctrl0_down_Decode_UOP_lane0;
      execute_ctrl1_up_Prediction_ALIGNED_JUMPED_lane0 <= execute_ctrl0_down_Prediction_ALIGNED_JUMPED_lane0;
      execute_ctrl1_up_Prediction_ALIGNED_JUMPED_PC_lane0 <= execute_ctrl0_down_Prediction_ALIGNED_JUMPED_PC_lane0;
      execute_ctrl1_up_Prediction_ALIGNED_SLICES_TAKEN_lane0 <= execute_ctrl0_down_Prediction_ALIGNED_SLICES_TAKEN_lane0;
      execute_ctrl1_up_Prediction_ALIGNED_SLICES_BRANCH_lane0 <= execute_ctrl0_down_Prediction_ALIGNED_SLICES_BRANCH_lane0;
      execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane0_0 <= execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane0_0;
      execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane0_1 <= execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane0_1;
      execute_ctrl1_up_Prediction_BRANCH_HISTORY_lane0 <= execute_ctrl0_down_Prediction_BRANCH_HISTORY_lane0;
      execute_ctrl1_up_Decode_INSTRUCTION_SLICE_COUNT_lane0 <= execute_ctrl0_down_Decode_INSTRUCTION_SLICE_COUNT_lane0;
      execute_ctrl1_up_PC_lane0 <= execute_ctrl0_down_PC_lane0;
      execute_ctrl1_up_TRAP_lane0 <= execute_ctrl0_down_TRAP_lane0;
      execute_ctrl1_up_Decode_UOP_ID_lane0 <= execute_ctrl0_down_Decode_UOP_ID_lane0;
      execute_ctrl1_up_RS1_PHYS_lane0 <= execute_ctrl0_down_RS1_PHYS_lane0;
      execute_ctrl1_up_RS2_PHYS_lane0 <= execute_ctrl0_down_RS2_PHYS_lane0;
      execute_ctrl1_up_RD_ENABLE_lane0 <= execute_ctrl0_down_RD_ENABLE_lane0;
      execute_ctrl1_up_RD_PHYS_lane0 <= execute_ctrl0_down_RD_PHYS_lane0;
      execute_ctrl1_up_COMPLETED_lane0 <= execute_ctrl0_down_COMPLETED_lane0;
      execute_ctrl1_up_AguPlugin_SIZE_lane0 <= execute_ctrl0_down_AguPlugin_SIZE_lane0;
    end
    if(execute_ctrl1_down_isReady) begin
      execute_ctrl2_up_Decode_UOP_lane0 <= execute_ctrl1_down_Decode_UOP_lane0;
      execute_ctrl2_up_Prediction_ALIGNED_JUMPED_lane0 <= execute_ctrl1_down_Prediction_ALIGNED_JUMPED_lane0;
      execute_ctrl2_up_Prediction_ALIGNED_JUMPED_PC_lane0 <= execute_ctrl1_down_Prediction_ALIGNED_JUMPED_PC_lane0;
      execute_ctrl2_up_Prediction_ALIGNED_SLICES_TAKEN_lane0 <= execute_ctrl1_down_Prediction_ALIGNED_SLICES_TAKEN_lane0;
      execute_ctrl2_up_Prediction_ALIGNED_SLICES_BRANCH_lane0 <= execute_ctrl1_down_Prediction_ALIGNED_SLICES_BRANCH_lane0;
      execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane0_0 <= execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane0_0;
      execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane0_1 <= execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane0_1;
      execute_ctrl2_up_Prediction_BRANCH_HISTORY_lane0 <= execute_ctrl1_down_Prediction_BRANCH_HISTORY_lane0;
      execute_ctrl2_up_Decode_INSTRUCTION_SLICE_COUNT_lane0 <= execute_ctrl1_down_Decode_INSTRUCTION_SLICE_COUNT_lane0;
      execute_ctrl2_up_PC_lane0 <= execute_ctrl1_down_PC_lane0;
      execute_ctrl2_up_TRAP_lane0 <= execute_ctrl1_down_TRAP_lane0;
      execute_ctrl2_up_Decode_UOP_ID_lane0 <= execute_ctrl1_down_Decode_UOP_ID_lane0;
      execute_ctrl2_up_RD_ENABLE_lane0 <= execute_ctrl1_down_RD_ENABLE_lane0;
      execute_ctrl2_up_RD_PHYS_lane0 <= execute_ctrl1_down_RD_PHYS_lane0;
      execute_ctrl2_up_COMPLETED_lane0 <= execute_ctrl1_down_COMPLETED_lane0;
      execute_ctrl2_up_AguPlugin_SIZE_lane0 <= execute_ctrl1_down_AguPlugin_SIZE_lane0;
      execute_ctrl2_up_early0_SrcPlugin_SRC1_lane0 <= execute_ctrl1_down_early0_SrcPlugin_SRC1_lane0;
      execute_ctrl2_up_integer_RS1_lane0 <= execute_ctrl1_down_integer_RS1_lane0;
      execute_ctrl2_up_early0_SrcPlugin_SRC2_lane0 <= execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0;
      execute_ctrl2_up_integer_RS2_lane0 <= execute_ctrl1_down_integer_RS2_lane0;
      execute_ctrl2_up_MAY_FLUSH_PRECISE_3_lane0 <= execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane0;
      execute_ctrl2_up_early0_IntAluPlugin_SEL_lane0 <= execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0;
      execute_ctrl2_up_early0_BarrelShifterPlugin_SEL_lane0 <= execute_ctrl1_down_early0_BarrelShifterPlugin_SEL_lane0;
      execute_ctrl2_up_early0_BranchPlugin_SEL_lane0 <= execute_ctrl1_down_early0_BranchPlugin_SEL_lane0;
      execute_ctrl2_up_early0_MulPlugin_SEL_lane0 <= execute_ctrl1_down_early0_MulPlugin_SEL_lane0;
      execute_ctrl2_up_early0_DivPlugin_SEL_lane0 <= execute_ctrl1_down_early0_DivPlugin_SEL_lane0;
      execute_ctrl2_up_early0_EnvPlugin_SEL_lane0 <= execute_ctrl1_down_early0_EnvPlugin_SEL_lane0;
      execute_ctrl2_up_MulPlugin_HIGH_lane0 <= execute_ctrl1_down_MulPlugin_HIGH_lane0;
      execute_ctrl2_up_CsrAccessPlugin_SEL_lane0 <= execute_ctrl1_down_CsrAccessPlugin_SEL_lane0;
      execute_ctrl2_up_AguPlugin_SEL_lane0 <= execute_ctrl1_down_AguPlugin_SEL_lane0;
      execute_ctrl2_up_LsuPlugin_logic_FENCE_lane0 <= execute_ctrl1_down_LsuPlugin_logic_FENCE_lane0;
      execute_ctrl2_up_lane0_integer_WriteBackPlugin_SEL_lane0 <= execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0;
      execute_ctrl2_up_COMPLETION_AT_2_lane0 <= execute_ctrl1_down_COMPLETION_AT_2_lane0;
      execute_ctrl2_up_COMPLETION_AT_4_lane0 <= execute_ctrl1_down_COMPLETION_AT_4_lane0;
      execute_ctrl2_up_COMPLETION_AT_3_lane0 <= execute_ctrl1_down_COMPLETION_AT_3_lane0;
      execute_ctrl2_up_lane0_logic_completions_onCtrl_0_ENABLE_lane0 <= execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0;
      execute_ctrl2_up_lane0_logic_completions_onCtrl_1_ENABLE_lane0 <= execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
      execute_ctrl2_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0 <= execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
      execute_ctrl2_up_early0_IntAluPlugin_ALU_ADD_SUB_lane0 <= execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0;
      execute_ctrl2_up_early0_IntAluPlugin_ALU_SLTX_lane0 <= execute_ctrl1_down_early0_IntAluPlugin_ALU_SLTX_lane0;
      execute_ctrl2_up_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0 <= execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
      execute_ctrl2_up_SrcStageables_REVERT_lane0 <= execute_ctrl1_down_SrcStageables_REVERT_lane0;
      execute_ctrl2_up_SrcStageables_ZERO_lane0 <= execute_ctrl1_down_SrcStageables_ZERO_lane0;
      execute_ctrl2_up_lane0_IntFormatPlugin_logic_SIGNED_lane0 <= execute_ctrl1_down_lane0_IntFormatPlugin_logic_SIGNED_lane0;
      execute_ctrl2_up_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0 <= execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
      execute_ctrl2_up_BYPASSED_AT_3_lane0 <= execute_ctrl1_down_BYPASSED_AT_3_lane0;
      execute_ctrl2_up_SrcStageables_UNSIGNED_lane0 <= execute_ctrl1_down_SrcStageables_UNSIGNED_lane0;
      execute_ctrl2_up_BarrelShifterPlugin_LEFT_lane0 <= execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0;
      execute_ctrl2_up_BarrelShifterPlugin_SIGNED_lane0 <= execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane0;
      execute_ctrl2_up_BarrelShifterPlugin_IS_W_lane0 <= execute_ctrl1_down_BarrelShifterPlugin_IS_W_lane0;
      execute_ctrl2_up_BarrelShifterPlugin_IS_W_RIGHT_lane0 <= execute_ctrl1_down_BarrelShifterPlugin_IS_W_RIGHT_lane0;
      execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane0 <= execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0;
      execute_ctrl2_up_RsUnsignedPlugin_RS1_SIGNED_lane0 <= execute_ctrl1_down_RsUnsignedPlugin_RS1_SIGNED_lane0;
      execute_ctrl2_up_RsUnsignedPlugin_RS2_SIGNED_lane0 <= execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0;
      execute_ctrl2_up_DivPlugin_REM_lane0 <= execute_ctrl1_down_DivPlugin_REM_lane0;
      execute_ctrl2_up_RsUnsignedPlugin_IS_W_lane0 <= execute_ctrl1_down_RsUnsignedPlugin_IS_W_lane0;
      execute_ctrl2_up_CsrAccessPlugin_CSR_IMM_lane0 <= execute_ctrl1_down_CsrAccessPlugin_CSR_IMM_lane0;
      execute_ctrl2_up_CsrAccessPlugin_CSR_MASK_lane0 <= execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0;
      execute_ctrl2_up_CsrAccessPlugin_CSR_CLEAR_lane0 <= execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0;
      execute_ctrl2_up_AguPlugin_LOAD_lane0 <= execute_ctrl1_down_AguPlugin_LOAD_lane0;
      execute_ctrl2_up_AguPlugin_STORE_lane0 <= execute_ctrl1_down_AguPlugin_STORE_lane0;
      execute_ctrl2_up_AguPlugin_ATOMIC_lane0 <= execute_ctrl1_down_AguPlugin_ATOMIC_lane0;
      execute_ctrl2_up_AguPlugin_FLOAT_lane0 <= execute_ctrl1_down_AguPlugin_FLOAT_lane0;
      execute_ctrl2_up_AguPlugin_CLEAN_lane0 <= execute_ctrl1_down_AguPlugin_CLEAN_lane0;
      execute_ctrl2_up_AguPlugin_INVALIDATE_lane0 <= execute_ctrl1_down_AguPlugin_INVALIDATE_lane0;
      execute_ctrl2_up_LsuPlugin_logic_LSU_PREFETCH_lane0 <= execute_ctrl1_down_LsuPlugin_logic_LSU_PREFETCH_lane0;
      execute_ctrl2_up_early0_EnvPlugin_OP_lane0 <= execute_ctrl1_down_early0_EnvPlugin_OP_lane0;
    end
    if(execute_ctrl2_down_isReady) begin
      execute_ctrl3_up_Decode_UOP_lane0 <= execute_ctrl2_down_Decode_UOP_lane0;
      execute_ctrl3_up_Prediction_BRANCH_HISTORY_lane0 <= execute_ctrl2_down_Prediction_BRANCH_HISTORY_lane0;
      execute_ctrl3_up_Decode_INSTRUCTION_SLICE_COUNT_lane0 <= execute_ctrl2_down_Decode_INSTRUCTION_SLICE_COUNT_lane0;
      execute_ctrl3_up_PC_lane0 <= execute_ctrl2_down_PC_lane0;
      execute_ctrl3_up_TRAP_lane0 <= execute_ctrl2_down_TRAP_lane0;
      execute_ctrl3_up_Decode_UOP_ID_lane0 <= execute_ctrl2_down_Decode_UOP_ID_lane0;
      execute_ctrl3_up_RD_ENABLE_lane0 <= execute_ctrl2_down_RD_ENABLE_lane0;
      execute_ctrl3_up_RD_PHYS_lane0 <= execute_ctrl2_down_RD_PHYS_lane0;
      execute_ctrl3_up_COMPLETED_lane0 <= execute_ctrl2_down_COMPLETED_lane0;
      execute_ctrl3_up_AguPlugin_SIZE_lane0 <= execute_ctrl2_down_AguPlugin_SIZE_lane0;
      execute_ctrl3_up_integer_RS2_lane0 <= execute_ctrl2_down_integer_RS2_lane0;
      execute_ctrl3_up_early0_MulPlugin_SEL_lane0 <= execute_ctrl2_down_early0_MulPlugin_SEL_lane0;
      execute_ctrl3_up_early0_DivPlugin_SEL_lane0 <= execute_ctrl2_down_early0_DivPlugin_SEL_lane0;
      execute_ctrl3_up_MulPlugin_HIGH_lane0 <= execute_ctrl2_down_MulPlugin_HIGH_lane0;
      execute_ctrl3_up_CsrAccessPlugin_SEL_lane0 <= execute_ctrl2_down_CsrAccessPlugin_SEL_lane0;
      execute_ctrl3_up_AguPlugin_SEL_lane0 <= execute_ctrl2_down_AguPlugin_SEL_lane0;
      execute_ctrl3_up_LsuPlugin_logic_FENCE_lane0 <= execute_ctrl2_down_LsuPlugin_logic_FENCE_lane0;
      execute_ctrl3_up_lane0_integer_WriteBackPlugin_SEL_lane0 <= execute_ctrl2_down_lane0_integer_WriteBackPlugin_SEL_lane0;
      execute_ctrl3_up_COMPLETION_AT_4_lane0 <= execute_ctrl2_down_COMPLETION_AT_4_lane0;
      execute_ctrl3_up_COMPLETION_AT_3_lane0 <= execute_ctrl2_down_COMPLETION_AT_3_lane0;
      execute_ctrl3_up_lane0_logic_completions_onCtrl_1_ENABLE_lane0 <= execute_ctrl2_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
      execute_ctrl3_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0 <= execute_ctrl2_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
      execute_ctrl3_up_lane0_IntFormatPlugin_logic_SIGNED_lane0 <= execute_ctrl2_down_lane0_IntFormatPlugin_logic_SIGNED_lane0;
      execute_ctrl3_up_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0 <= execute_ctrl2_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
      execute_ctrl3_up_AguPlugin_LOAD_lane0 <= execute_ctrl2_down_AguPlugin_LOAD_lane0;
      execute_ctrl3_up_AguPlugin_STORE_lane0 <= execute_ctrl2_down_AguPlugin_STORE_lane0;
      execute_ctrl3_up_AguPlugin_ATOMIC_lane0 <= execute_ctrl2_down_AguPlugin_ATOMIC_lane0;
      execute_ctrl3_up_AguPlugin_FLOAT_lane0 <= execute_ctrl2_down_AguPlugin_FLOAT_lane0;
      execute_ctrl3_up_LsuPlugin_logic_LSU_PREFETCH_lane0 <= execute_ctrl2_down_LsuPlugin_logic_LSU_PREFETCH_lane0;
      execute_ctrl3_up_LsuL1Plugin_logic_FREEZE_HAZARD_lane0 <= execute_ctrl2_down_LsuL1Plugin_logic_FREEZE_HAZARD_lane0;
      execute_ctrl3_up_COMMIT_lane0 <= execute_ctrl2_down_COMMIT_lane0;
      execute_ctrl3_up_early0_SrcPlugin_ADD_SUB_lane0 <= execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0;
      execute_ctrl3_up_LsuL1_MIXED_ADDRESS_lane0 <= execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0;
      execute_ctrl3_up_LsuL1Plugin_logic_BANK_BUSY_lane0 <= execute_ctrl2_down_LsuL1Plugin_logic_BANK_BUSY_lane0;
      execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_VALID_lane0 <= execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_VALID_lane0;
      execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_ADDRESS_lane0 <= execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_ADDRESS_lane0;
      execute_ctrl3_up_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALID_lane0 <= execute_ctrl2_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALID_lane0;
      execute_ctrl3_up_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_plru_0 <= execute_ctrl2_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_plru_0;
      execute_ctrl3_up_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_dirty <= execute_ctrl2_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_dirty;
      execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0 <= execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0;
      execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0 <= execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0;
      execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_0_lane0 <= execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_0_lane0;
      execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_1_lane0 <= execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_1_lane0;
      execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_2_lane0 <= execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_2_lane0;
      execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_3_lane0 <= execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_3_lane0;
      execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_4_lane0 <= execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_4_lane0;
      execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_5_lane0 <= execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_5_lane0;
      execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_6_lane0 <= execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_6_lane0;
      execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_7_lane0 <= execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_7_lane0;
      execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_8_lane0 <= execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_8_lane0;
      execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_9_lane0 <= execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_9_lane0;
      execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_10_lane0 <= execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_10_lane0;
      execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_11_lane0 <= execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_11_lane0;
      execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_12_lane0 <= execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_12_lane0;
      execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_13_lane0 <= execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_13_lane0;
      execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_14_lane0 <= execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_14_lane0;
      execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_15_lane0 <= execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_15_lane0;
      execute_ctrl3_up_DivPlugin_DIV_RESULT_lane0 <= execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0;
      execute_ctrl3_up_LsuPlugin_logic_FORCE_PHYSICAL_lane0 <= execute_ctrl2_down_LsuPlugin_logic_FORCE_PHYSICAL_lane0;
      execute_ctrl3_up_LsuPlugin_logic_FROM_ACCESS_lane0 <= execute_ctrl2_down_LsuPlugin_logic_FROM_ACCESS_lane0;
      execute_ctrl3_up_LsuL1_MASK_lane0 <= execute_ctrl2_down_LsuL1_MASK_lane0;
      execute_ctrl3_up_LsuL1_SIZE_lane0 <= execute_ctrl2_down_LsuL1_SIZE_lane0;
      execute_ctrl3_up_LsuL1_LOAD_lane0 <= execute_ctrl2_down_LsuL1_LOAD_lane0;
      execute_ctrl3_up_LsuL1_ATOMIC_lane0 <= execute_ctrl2_down_LsuL1_ATOMIC_lane0;
      execute_ctrl3_up_LsuL1_STORE_lane0 <= execute_ctrl2_down_LsuL1_STORE_lane0;
      execute_ctrl3_up_LsuL1_CLEAN_lane0 <= execute_ctrl2_down_LsuL1_CLEAN_lane0;
      execute_ctrl3_up_LsuL1_INVALID_lane0 <= execute_ctrl2_down_LsuL1_INVALID_lane0;
      execute_ctrl3_up_LsuL1_PREFETCH_lane0 <= execute_ctrl2_down_LsuL1_PREFETCH_lane0;
      execute_ctrl3_up_LsuL1_FLUSH_lane0 <= execute_ctrl2_down_LsuL1_FLUSH_lane0;
      execute_ctrl3_up_Decode_STORE_ID_lane0 <= execute_ctrl2_down_Decode_STORE_ID_lane0;
      execute_ctrl3_up_LsuPlugin_logic_FROM_LSU_lane0 <= execute_ctrl2_down_LsuPlugin_logic_FROM_LSU_lane0;
      execute_ctrl3_up_LsuPlugin_logic_FROM_PREFETCH_lane0 <= execute_ctrl2_down_LsuPlugin_logic_FROM_PREFETCH_lane0;
      execute_ctrl3_up_LsuPlugin_logic_pmpPort_logic_onEntries_0_PERM_OK_lane0 <= execute_ctrl2_down_LsuPlugin_logic_pmpPort_logic_onEntries_0_PERM_OK_lane0;
      execute_ctrl3_up_LsuPlugin_logic_pmpPort_logic_onEntries_1_PERM_OK_lane0 <= execute_ctrl2_down_LsuPlugin_logic_pmpPort_logic_onEntries_1_PERM_OK_lane0;
      execute_ctrl3_up_LsuPlugin_logic_pmpPort_logic_onEntries_2_PERM_OK_lane0 <= execute_ctrl2_down_LsuPlugin_logic_pmpPort_logic_onEntries_2_PERM_OK_lane0;
      execute_ctrl3_up_LsuPlugin_logic_pmpPort_logic_onEntries_3_PERM_OK_lane0 <= execute_ctrl2_down_LsuPlugin_logic_pmpPort_logic_onEntries_3_PERM_OK_lane0;
      execute_ctrl3_up_LsuPlugin_logic_pmpPort_logic_NEED_HIT_lane0 <= execute_ctrl2_down_LsuPlugin_logic_pmpPort_logic_NEED_HIT_lane0;
      execute_ctrl3_up_lane0_integer_WriteBackPlugin_logic_DATA_lane0 <= execute_ctrl2_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
      execute_ctrl3_up_MMU_L0_ENTRIES_lane0_0_valid <= execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_valid;
      execute_ctrl3_up_MMU_L0_ENTRIES_lane0_0_virtualAddress <= execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_virtualAddress;
      execute_ctrl3_up_MMU_L0_ENTRIES_lane0_0_physicalAddress <= execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_physicalAddress;
      execute_ctrl3_up_MMU_L0_ENTRIES_lane0_0_allowRead <= execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_allowRead;
      execute_ctrl3_up_MMU_L0_ENTRIES_lane0_0_allowWrite <= execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_allowWrite;
      execute_ctrl3_up_MMU_L0_ENTRIES_lane0_0_allowExecute <= execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_allowExecute;
      execute_ctrl3_up_MMU_L0_ENTRIES_lane0_0_allowUser <= execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_allowUser;
      execute_ctrl3_up_MMU_L0_ENTRIES_lane0_1_valid <= execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_valid;
      execute_ctrl3_up_MMU_L0_ENTRIES_lane0_1_virtualAddress <= execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_virtualAddress;
      execute_ctrl3_up_MMU_L0_ENTRIES_lane0_1_physicalAddress <= execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_physicalAddress;
      execute_ctrl3_up_MMU_L0_ENTRIES_lane0_1_allowRead <= execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_allowRead;
      execute_ctrl3_up_MMU_L0_ENTRIES_lane0_1_allowWrite <= execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_allowWrite;
      execute_ctrl3_up_MMU_L0_ENTRIES_lane0_1_allowExecute <= execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_allowExecute;
      execute_ctrl3_up_MMU_L0_ENTRIES_lane0_1_allowUser <= execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_allowUser;
      execute_ctrl3_up_MMU_L0_ENTRIES_lane0_2_valid <= execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_valid;
      execute_ctrl3_up_MMU_L0_ENTRIES_lane0_2_virtualAddress <= execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_virtualAddress;
      execute_ctrl3_up_MMU_L0_ENTRIES_lane0_2_physicalAddress <= execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_physicalAddress;
      execute_ctrl3_up_MMU_L0_ENTRIES_lane0_2_allowRead <= execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_allowRead;
      execute_ctrl3_up_MMU_L0_ENTRIES_lane0_2_allowWrite <= execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_allowWrite;
      execute_ctrl3_up_MMU_L0_ENTRIES_lane0_2_allowExecute <= execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_allowExecute;
      execute_ctrl3_up_MMU_L0_ENTRIES_lane0_2_allowUser <= execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_allowUser;
      execute_ctrl3_up_MMU_L0_HITS_PRE_VALID_lane0 <= execute_ctrl2_down_MMU_L0_HITS_PRE_VALID_lane0;
      execute_ctrl3_up_MMU_L1_ENTRIES_lane0_0_valid <= execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_valid;
      execute_ctrl3_up_MMU_L1_ENTRIES_lane0_0_virtualAddress <= execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_virtualAddress;
      execute_ctrl3_up_MMU_L1_ENTRIES_lane0_0_physicalAddress <= execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_physicalAddress;
      execute_ctrl3_up_MMU_L1_ENTRIES_lane0_0_allowRead <= execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_allowRead;
      execute_ctrl3_up_MMU_L1_ENTRIES_lane0_0_allowWrite <= execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_allowWrite;
      execute_ctrl3_up_MMU_L1_ENTRIES_lane0_0_allowExecute <= execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_allowExecute;
      execute_ctrl3_up_MMU_L1_ENTRIES_lane0_0_allowUser <= execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_allowUser;
      execute_ctrl3_up_MMU_L1_HITS_PRE_VALID_lane0 <= execute_ctrl2_down_MMU_L1_HITS_PRE_VALID_lane0;
    end
    if(execute_ctrl3_down_isReady) begin
      execute_ctrl4_up_Decode_UOP_lane0 <= execute_ctrl3_down_Decode_UOP_lane0;
      execute_ctrl4_up_Prediction_BRANCH_HISTORY_lane0 <= execute_ctrl3_down_Prediction_BRANCH_HISTORY_lane0;
      execute_ctrl4_up_Decode_INSTRUCTION_SLICE_COUNT_lane0 <= execute_ctrl3_down_Decode_INSTRUCTION_SLICE_COUNT_lane0;
      execute_ctrl4_up_PC_lane0 <= execute_ctrl3_down_PC_lane0;
      execute_ctrl4_up_TRAP_lane0 <= execute_ctrl3_down_TRAP_lane0;
      execute_ctrl4_up_Decode_UOP_ID_lane0 <= execute_ctrl3_down_Decode_UOP_ID_lane0;
      execute_ctrl4_up_RD_ENABLE_lane0 <= execute_ctrl3_down_RD_ENABLE_lane0;
      execute_ctrl4_up_RD_PHYS_lane0 <= execute_ctrl3_down_RD_PHYS_lane0;
      execute_ctrl4_up_COMPLETED_lane0 <= execute_ctrl3_down_COMPLETED_lane0;
      execute_ctrl4_up_AguPlugin_SIZE_lane0 <= execute_ctrl3_down_AguPlugin_SIZE_lane0;
      execute_ctrl4_up_integer_RS2_lane0 <= execute_ctrl3_down_integer_RS2_lane0;
      execute_ctrl4_up_early0_MulPlugin_SEL_lane0 <= execute_ctrl3_down_early0_MulPlugin_SEL_lane0;
      execute_ctrl4_up_MulPlugin_HIGH_lane0 <= execute_ctrl3_down_MulPlugin_HIGH_lane0;
      execute_ctrl4_up_AguPlugin_SEL_lane0 <= execute_ctrl3_down_AguPlugin_SEL_lane0;
      execute_ctrl4_up_LsuPlugin_logic_FENCE_lane0 <= execute_ctrl3_down_LsuPlugin_logic_FENCE_lane0;
      execute_ctrl4_up_lane0_integer_WriteBackPlugin_SEL_lane0 <= execute_ctrl3_down_lane0_integer_WriteBackPlugin_SEL_lane0;
      execute_ctrl4_up_COMPLETION_AT_4_lane0 <= execute_ctrl3_down_COMPLETION_AT_4_lane0;
      execute_ctrl4_up_lane0_logic_completions_onCtrl_1_ENABLE_lane0 <= execute_ctrl3_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
      execute_ctrl4_up_lane0_IntFormatPlugin_logic_SIGNED_lane0 <= execute_ctrl3_down_lane0_IntFormatPlugin_logic_SIGNED_lane0;
      execute_ctrl4_up_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0 <= execute_ctrl3_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
      execute_ctrl4_up_AguPlugin_LOAD_lane0 <= execute_ctrl3_down_AguPlugin_LOAD_lane0;
      execute_ctrl4_up_AguPlugin_STORE_lane0 <= execute_ctrl3_down_AguPlugin_STORE_lane0;
      execute_ctrl4_up_AguPlugin_ATOMIC_lane0 <= execute_ctrl3_down_AguPlugin_ATOMIC_lane0;
      execute_ctrl4_up_AguPlugin_FLOAT_lane0 <= execute_ctrl3_down_AguPlugin_FLOAT_lane0;
      execute_ctrl4_up_LsuPlugin_logic_LSU_PREFETCH_lane0 <= execute_ctrl3_down_LsuPlugin_logic_LSU_PREFETCH_lane0;
      execute_ctrl4_up_LsuL1Plugin_logic_FREEZE_HAZARD_lane0 <= execute_ctrl3_down_LsuL1Plugin_logic_FREEZE_HAZARD_lane0;
      execute_ctrl4_up_COMMIT_lane0 <= execute_ctrl3_down_COMMIT_lane0;
      execute_ctrl4_up_LsuL1_MIXED_ADDRESS_lane0 <= execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0;
      execute_ctrl4_up_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0 <= execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0;
      execute_ctrl4_up_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0 <= execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0;
      execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_0_lane0 <= execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_0_lane0;
      execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_1_lane0 <= execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_1_lane0;
      execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_2_lane0 <= execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_2_lane0;
      execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_3_lane0 <= execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_3_lane0;
      execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_4_lane0 <= execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_4_lane0;
      execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_5_lane0 <= execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_5_lane0;
      execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_6_lane0 <= execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_6_lane0;
      execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_7_lane0 <= execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_7_lane0;
      execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_8_lane0 <= execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_8_lane0;
      execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_9_lane0 <= execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_9_lane0;
      execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_10_lane0 <= execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_10_lane0;
      execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_11_lane0 <= execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_11_lane0;
      execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_12_lane0 <= execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_12_lane0;
      execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_13_lane0 <= execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_13_lane0;
      execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_14_lane0 <= execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_14_lane0;
      execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_15_lane0 <= execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_15_lane0;
      execute_ctrl4_up_LsuPlugin_logic_FROM_ACCESS_lane0 <= execute_ctrl3_down_LsuPlugin_logic_FROM_ACCESS_lane0;
      execute_ctrl4_up_LsuL1_MASK_lane0 <= execute_ctrl3_down_LsuL1_MASK_lane0;
      execute_ctrl4_up_LsuL1_SIZE_lane0 <= execute_ctrl3_down_LsuL1_SIZE_lane0;
      execute_ctrl4_up_LsuL1_LOAD_lane0 <= execute_ctrl3_down_LsuL1_LOAD_lane0;
      execute_ctrl4_up_LsuL1_ATOMIC_lane0 <= execute_ctrl3_down_LsuL1_ATOMIC_lane0;
      execute_ctrl4_up_LsuL1_STORE_lane0 <= execute_ctrl3_down_LsuL1_STORE_lane0;
      execute_ctrl4_up_LsuL1_CLEAN_lane0 <= execute_ctrl3_down_LsuL1_CLEAN_lane0;
      execute_ctrl4_up_LsuL1_INVALID_lane0 <= execute_ctrl3_down_LsuL1_INVALID_lane0;
      execute_ctrl4_up_LsuL1_PREFETCH_lane0 <= execute_ctrl3_down_LsuL1_PREFETCH_lane0;
      execute_ctrl4_up_LsuL1_FLUSH_lane0 <= execute_ctrl3_down_LsuL1_FLUSH_lane0;
      execute_ctrl4_up_Decode_STORE_ID_lane0 <= execute_ctrl3_down_Decode_STORE_ID_lane0;
      execute_ctrl4_up_LsuPlugin_logic_FROM_LSU_lane0 <= execute_ctrl3_down_LsuPlugin_logic_FROM_LSU_lane0;
      execute_ctrl4_up_LsuPlugin_logic_FROM_PREFETCH_lane0 <= execute_ctrl3_down_LsuPlugin_logic_FROM_PREFETCH_lane0;
      execute_ctrl4_up_LsuPlugin_logic_pmpPort_logic_onEntries_0_PERM_OK_lane0 <= execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_0_PERM_OK_lane0;
      execute_ctrl4_up_LsuPlugin_logic_pmpPort_logic_onEntries_1_PERM_OK_lane0 <= execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_1_PERM_OK_lane0;
      execute_ctrl4_up_LsuPlugin_logic_pmpPort_logic_onEntries_2_PERM_OK_lane0 <= execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_2_PERM_OK_lane0;
      execute_ctrl4_up_LsuPlugin_logic_pmpPort_logic_onEntries_3_PERM_OK_lane0 <= execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_3_PERM_OK_lane0;
      execute_ctrl4_up_LsuPlugin_logic_pmpPort_logic_NEED_HIT_lane0 <= execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_NEED_HIT_lane0;
      execute_ctrl4_up_lane0_integer_WriteBackPlugin_logic_DATA_lane0 <= execute_ctrl3_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
      execute_ctrl4_up_LsuL1Plugin_logic_SHARED_lane0_plru_0 <= execute_ctrl3_down_LsuL1Plugin_logic_SHARED_lane0_plru_0;
      execute_ctrl4_up_LsuL1Plugin_logic_SHARED_lane0_dirty <= execute_ctrl3_down_LsuL1Plugin_logic_SHARED_lane0_dirty;
      execute_ctrl4_up_LsuL1Plugin_logic_BANK_BUSY_REMAPPED_lane0 <= execute_ctrl3_down_LsuL1Plugin_logic_BANK_BUSY_REMAPPED_lane0;
      execute_ctrl4_up_LsuL1Plugin_logic_BANKS_MUXES_lane0_0 <= execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0;
      execute_ctrl4_up_LsuL1Plugin_logic_BANKS_MUXES_lane0_1 <= execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1;
      execute_ctrl4_up_LsuL1Plugin_logic_WRITE_TO_READ_HAZARDS_lane0 <= execute_ctrl3_down_LsuL1Plugin_logic_WRITE_TO_READ_HAZARDS_lane0;
      execute_ctrl4_up_LsuL1_PHYSICAL_ADDRESS_lane0 <= execute_ctrl3_down_LsuL1_PHYSICAL_ADDRESS_lane0;
      execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_loaded <= execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_loaded;
      execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_address <= execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_address;
      execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault <= execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault;
      execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_loaded <= execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_loaded;
      execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_address <= execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_address;
      execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault <= execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault;
      execute_ctrl4_up_LsuL1Plugin_logic_WAYS_HITS_lane0 <= execute_ctrl3_down_LsuL1Plugin_logic_WAYS_HITS_lane0;
      execute_ctrl4_up_early0_MulPlugin_logic_steps_0_adders_0_lane0 <= execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0;
      execute_ctrl4_up_early0_MulPlugin_logic_steps_0_adders_1_lane0 <= execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0;
      execute_ctrl4_up_early0_MulPlugin_logic_steps_0_adders_2_lane0 <= execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0;
      execute_ctrl4_up_LsuPlugin_logic_onTrigger_HIT_lane0 <= execute_ctrl3_down_LsuPlugin_logic_onTrigger_HIT_lane0;
      execute_ctrl4_up_MMU_TRANSLATED_lane0 <= execute_ctrl3_down_MMU_TRANSLATED_lane0;
      execute_ctrl4_up_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0 <= execute_ctrl3_down_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0;
      execute_ctrl4_up_LsuPlugin_logic_preCtrl_IS_AMO_lane0 <= execute_ctrl3_down_LsuPlugin_logic_preCtrl_IS_AMO_lane0;
      execute_ctrl4_up_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault <= execute_ctrl3_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault;
      execute_ctrl4_up_LsuPlugin_logic_onPma_CACHED_RSP_lane0_io <= execute_ctrl3_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_io;
      execute_ctrl4_up_LsuPlugin_logic_onPma_IO_RSP_lane0_fault <= execute_ctrl3_down_LsuPlugin_logic_onPma_IO_RSP_lane0_fault;
      execute_ctrl4_up_LsuPlugin_logic_onPma_IO_RSP_lane0_io <= execute_ctrl3_down_LsuPlugin_logic_onPma_IO_RSP_lane0_io;
      execute_ctrl4_up_LsuPlugin_logic_onPma_IO_lane0 <= execute_ctrl3_down_LsuPlugin_logic_onPma_IO_lane0;
      execute_ctrl4_up_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0 <= execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0;
      execute_ctrl4_up_LsuPlugin_logic_MMU_PAGE_FAULT_lane0 <= execute_ctrl3_down_LsuPlugin_logic_MMU_PAGE_FAULT_lane0;
      execute_ctrl4_up_LsuPlugin_logic_MMU_FAILURE_lane0 <= execute_ctrl3_down_LsuPlugin_logic_MMU_FAILURE_lane0;
      execute_ctrl4_up_MMU_ACCESS_FAULT_lane0 <= execute_ctrl3_down_MMU_ACCESS_FAULT_lane0;
      execute_ctrl4_up_MMU_REFILL_lane0 <= execute_ctrl3_down_MMU_REFILL_lane0;
      execute_ctrl4_up_MMU_HAZARD_lane0 <= execute_ctrl3_down_MMU_HAZARD_lane0;
      execute_ctrl4_up_LsuPlugin_logic_pmpPort_logic_onEntries_0_napot_HIT_lane0 <= execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_0_napot_HIT_lane0;
      execute_ctrl4_up_LsuPlugin_logic_pmpPort_logic_onEntries_0_tor_BIGGER_lane0 <= execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_0_tor_BIGGER_lane0;
      execute_ctrl4_up_LsuPlugin_logic_pmpPort_logic_onEntries_1_napot_HIT_lane0 <= execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_1_napot_HIT_lane0;
      execute_ctrl4_up_LsuPlugin_logic_pmpPort_logic_onEntries_1_tor_BIGGER_lane0 <= execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_1_tor_BIGGER_lane0;
      execute_ctrl4_up_LsuPlugin_logic_pmpPort_logic_onEntries_2_napot_HIT_lane0 <= execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_2_napot_HIT_lane0;
      execute_ctrl4_up_LsuPlugin_logic_pmpPort_logic_onEntries_2_tor_BIGGER_lane0 <= execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_2_tor_BIGGER_lane0;
      execute_ctrl4_up_LsuPlugin_logic_pmpPort_logic_onEntries_3_napot_HIT_lane0 <= execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_3_napot_HIT_lane0;
      execute_ctrl4_up_LsuPlugin_logic_pmpPort_logic_onEntries_3_tor_BIGGER_lane0 <= execute_ctrl3_down_LsuPlugin_logic_pmpPort_logic_onEntries_3_tor_BIGGER_lane0;
      execute_ctrl4_up_MMU_BYPASS_TRANSLATION_lane0 <= execute_ctrl3_down_MMU_BYPASS_TRANSLATION_lane0;
    end
    if(execute_ctrl4_down_isReady) begin
      execute_ctrl5_up_RD_ENABLE_lane0 <= execute_ctrl4_down_RD_ENABLE_lane0;
      execute_ctrl5_up_RD_PHYS_lane0 <= execute_ctrl4_down_RD_PHYS_lane0;
      execute_ctrl5_up_COMMIT_lane0 <= execute_ctrl4_down_COMMIT_lane0;
      execute_ctrl5_up_lane0_integer_WriteBackPlugin_logic_DATA_lane0 <= execute_ctrl4_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
    end
    case(LsuPlugin_logic_flusher_stateReg)
      LsuPlugin_logic_flusher_CMD : begin
        if(when_LsuPlugin_l368) begin
          LsuPlugin_logic_flusher_waiter <= LsuL1_WRITEBACK_BUSY;
        end
      end
      LsuPlugin_logic_flusher_COMPLETION : begin
        LsuPlugin_logic_flusher_waiter <= (LsuPlugin_logic_flusher_waiter & LsuL1_WRITEBACK_BUSY);
      end
      default : begin
        LsuPlugin_logic_flusher_cmdCounter <= 7'h0;
      end
    endcase
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
        TrapPlugin_logic_harts_0_trap_fsm_triggerEbreakReg <= TrapPlugin_logic_harts_0_trap_fsm_triggerEbreak;
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_WAIT : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
        if(TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_valid) begin
          if(when_TrapPlugin_l555) begin
            TrapPlugin_logic_harts_0_trap_pending_state_exception <= 1'b1;
            case(switch_TrapPlugin_l557)
              3'b110 : begin
                TrapPlugin_logic_harts_0_trap_pending_state_code <= 4'b0001;
              end
              3'b100 : begin
                TrapPlugin_logic_harts_0_trap_pending_state_code <= 4'b0101;
              end
              3'b101 : begin
                TrapPlugin_logic_harts_0_trap_pending_state_code <= 4'b0111;
              end
              3'b010 : begin
                TrapPlugin_logic_harts_0_trap_pending_state_code <= 4'b1100;
              end
              3'b000 : begin
                TrapPlugin_logic_harts_0_trap_pending_state_code <= 4'b1101;
              end
              3'b001 : begin
                TrapPlugin_logic_harts_0_trap_pending_state_code <= 4'b1111;
              end
              default : begin
              end
            endcase
          end
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
        if(MmuPlugin_logic_refill_arbiter_io_output_valid) begin
          MmuPlugin_logic_refill_portOhReg <= MmuPlugin_logic_refill_arbiter_io_chosenOH;
          MmuPlugin_logic_refill_storageOhReg <= (2'b01 <<< MmuPlugin_logic_refill_arbiter_io_output_payload_storageId);
          MmuPlugin_logic_refill_storageEnable <= MmuPlugin_logic_refill_arbiter_io_output_payload_storageEnable;
          MmuPlugin_logic_refill_virtual <= MmuPlugin_logic_refill_arbiter_io_output_payload_address;
          MmuPlugin_logic_refill_load_address <= _zz_MmuPlugin_logic_refill_load_address[31:0];
        end
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_CMD_2 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(!when_MmuPlugin_l534) begin
              MmuPlugin_logic_refill_load_address <= MmuPlugin_logic_refill_load_nextLevelBase;
              MmuPlugin_logic_refill_load_address[11 : 3] <= MmuPlugin_logic_refill_virtual[20 : 12];
            end
          end
        end
      end
      MmuPlugin_logic_refill_RSP_2 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(!when_MmuPlugin_l534_1) begin
              MmuPlugin_logic_refill_load_address <= MmuPlugin_logic_refill_load_nextLevelBase;
              MmuPlugin_logic_refill_load_address[11 : 3] <= MmuPlugin_logic_refill_virtual[29 : 21];
            end
          end
        end
      end
      MmuPlugin_logic_refill_DONE_0 : begin
      end
      MmuPlugin_logic_refill_DONE_1 : begin
      end
      MmuPlugin_logic_refill_DONE_2 : begin
      end
      default : begin
      end
    endcase
    case(PerformanceCounterPlugin_logic_fsm_stateReg)
      PerformanceCounterPlugin_logic_fsm_IDLE : begin
        PerformanceCounterPlugin_logic_fsm_cmd_oh <= {(PerformanceCounterPlugin_logic_fsm_idleCsrAddress == 2'b10),(PerformanceCounterPlugin_logic_fsm_idleCsrAddress == 2'b00)};
        if(!PerformanceCounterPlugin_logic_fsm_csrWriteCmd_valid) begin
          if(PerformanceCounterPlugin_logic_fsm_flusherCmd_valid) begin
            PerformanceCounterPlugin_logic_fsm_cmd_flusher <= 1'b1;
            PerformanceCounterPlugin_logic_fsm_cmd_oh <= PerformanceCounterPlugin_logic_fsm_flusherCmd_payload_oh;
          end else begin
            if(PerformanceCounterPlugin_logic_fsm_csrReadCmd_valid) begin
              PerformanceCounterPlugin_logic_fsm_cmd_flusher <= 1'b0;
            end
          end
        end
        PerformanceCounterPlugin_logic_fsm_carry <= 1'b0;
      end
      PerformanceCounterPlugin_logic_fsm_READ_LOW : begin
        PerformanceCounterPlugin_logic_fsm_ramReaded <= PerformanceCounterPlugin_logic_readPort_data;
        PerformanceCounterPlugin_logic_fsm_counterReaded <= ((_zz_PerformanceCounterPlugin_logic_fsm_cmd_address ? PerformanceCounterPlugin_logic_counters_cycle_value : 8'h0) | (_zz_PerformanceCounterPlugin_logic_fsm_cmd_address_1 ? PerformanceCounterPlugin_logic_counters_instret_value : 8'h0));
      end
      PerformanceCounterPlugin_logic_fsm_CALC_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_CSR_WRITE : begin
      end
      default : begin
      end
    endcase
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_READ : begin
        CsrAccessPlugin_logic_fsm_interface_aluInput <= CsrAccessPlugin_bus_read_toWriteBits;
        CsrAccessPlugin_logic_fsm_interface_csrValue <= CsrAccessPlugin_logic_fsm_readLogic_csrValue;
      end
      CsrAccessPlugin_logic_fsm_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_COMPLETION : begin
      end
      default : begin
        REG_CSR_768 <= COMB_CSR_768;
        REG_CSR_256 <= COMB_CSR_256;
        REG_CSR_384 <= COMB_CSR_384;
        REG_CSR_944 <= COMB_CSR_944;
        REG_CSR_928 <= COMB_CSR_928;
        REG_CSR_945 <= COMB_CSR_945;
        REG_CSR_946 <= COMB_CSR_946;
        REG_CSR_947 <= COMB_CSR_947;
        REG_CSR_PmpPlugin_logic_allFilter <= COMB_CSR_PmpPlugin_logic_allFilter;
        REG_CSR_794 <= COMB_CSR_794;
        REG_CSR_1952 <= COMB_CSR_1952;
        REG_CSR_1953 <= COMB_CSR_1953;
        REG_CSR_1954 <= COMB_CSR_1954;
        REG_CSR_3857 <= COMB_CSR_3857;
        REG_CSR_3858 <= COMB_CSR_3858;
        REG_CSR_3859 <= COMB_CSR_3859;
        REG_CSR_3860 <= COMB_CSR_3860;
        REG_CSR_769 <= COMB_CSR_769;
        REG_CSR_834 <= COMB_CSR_834;
        REG_CSR_836 <= COMB_CSR_836;
        REG_CSR_772 <= COMB_CSR_772;
        REG_CSR_770 <= COMB_CSR_770;
        REG_CSR_771 <= COMB_CSR_771;
        REG_CSR_4016 <= COMB_CSR_4016;
        REG_CSR_774 <= COMB_CSR_774;
        REG_CSR_322 <= COMB_CSR_322;
        REG_CSR_778 <= COMB_CSR_778;
        REG_CSR_260 <= COMB_CSR_260;
        REG_CSR_324 <= COMB_CSR_324;
        REG_CSR_3504 <= COMB_CSR_3504;
        REG_CSR_3073 <= COMB_CSR_3073;
        REG_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_tvecFilter <= COMB_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_tvecFilter;
        REG_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_epcFilter <= COMB_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_epcFilter;
        REG_CSR_262 <= COMB_CSR_262;
        REG_CSR_800 <= COMB_CSR_800;
        REG_CSR_UNAMED_0 <= COMB_CSR_UNAMED_1;
        REG_CSR_266 <= COMB_CSR_266;
        REG_CSR_CsrRamPlugin_csrMapper_selFilter <= COMB_CSR_CsrRamPlugin_csrMapper_selFilter;
        REG_CSR_PerformanceCounterPlugin_logic_csrFilter <= COMB_CSR_PerformanceCounterPlugin_logic_csrFilter;
        REG_CSR_CsrAccessPlugin_logic_trapNextOnWriteFilter <= COMB_CSR_CsrAccessPlugin_logic_trapNextOnWriteFilter;
      end
    endcase
  end


endmodule

module RegFileMem (
  input  wire          io_writes_0_valid,
  input  wire [4:0]    io_writes_0_address,
  input  wire [63:0]   io_writes_0_data,
  input  wire [15:0]   io_writes_0_uopId,
  input  wire          io_reads_0_valid,
  input  wire [4:0]    io_reads_0_address,
  output wire [63:0]   io_reads_0_data,
  input  wire          io_reads_1_valid,
  input  wire [4:0]    io_reads_1_address,
  output wire [63:0]   io_reads_1_data,
  input  wire          clk,
  input  wire          reset
);

  reg        [63:0]   asMem_ram_spinal_port1;
  reg        [63:0]   asMem_ram_spinal_port2;
  reg                 _zz_1;
  wire                conv_writes_0_valid;
  wire       [4:0]    conv_writes_0_payload_address;
  wire       [63:0]   conv_writes_0_payload_data;
  wire                conv_read_0_cmd_valid;
  wire       [4:0]    conv_read_0_cmd_payload;
  wire       [63:0]   conv_read_0_rsp;
  wire                conv_read_1_cmd_valid;
  wire       [4:0]    conv_read_1_cmd_payload;
  wire       [63:0]   conv_read_1_rsp;
  wire                asMem_writes_0_port_valid;
  wire       [4:0]    asMem_writes_0_port_payload_address;
  wire       [63:0]   asMem_writes_0_port_payload_data;
  wire                asMem_reads_0_sync_port_cmd_valid;
  wire       [4:0]    asMem_reads_0_sync_port_cmd_payload;
  wire       [63:0]   asMem_reads_0_sync_port_rsp;
  wire                asMem_reads_1_sync_port_cmd_valid;
  wire       [4:0]    asMem_reads_1_sync_port_cmd_payload;
  wire       [63:0]   asMem_reads_1_sync_port_rsp;
  reg [63:0] asMem_ram [0:31] /* verilator public */ ;

  always @(posedge clk) begin
    if(_zz_1) begin
      asMem_ram[asMem_writes_0_port_payload_address] <= asMem_writes_0_port_payload_data;
    end
  end

  always @(posedge clk) begin
    if(asMem_reads_0_sync_port_cmd_valid) begin
      asMem_ram_spinal_port1 <= asMem_ram[asMem_reads_0_sync_port_cmd_payload];
    end
  end

  always @(posedge clk) begin
    if(asMem_reads_1_sync_port_cmd_valid) begin
      asMem_ram_spinal_port2 <= asMem_ram[asMem_reads_1_sync_port_cmd_payload];
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(asMem_writes_0_port_valid) begin
      _zz_1 = 1'b1;
    end
  end

  assign conv_writes_0_valid = io_writes_0_valid;
  assign conv_writes_0_payload_address = io_writes_0_address;
  assign conv_writes_0_payload_data = io_writes_0_data;
  assign conv_read_0_cmd_valid = io_reads_0_valid;
  assign conv_read_0_cmd_payload = io_reads_0_address;
  assign io_reads_0_data = conv_read_0_rsp;
  assign conv_read_1_cmd_valid = io_reads_1_valid;
  assign conv_read_1_cmd_payload = io_reads_1_address;
  assign io_reads_1_data = conv_read_1_rsp;
  assign asMem_writes_0_port_valid = conv_writes_0_valid;
  assign asMem_writes_0_port_payload_address = conv_writes_0_payload_address;
  assign asMem_writes_0_port_payload_data = conv_writes_0_payload_data;
  assign asMem_reads_0_sync_port_rsp = asMem_ram_spinal_port1;
  assign asMem_reads_0_sync_port_cmd_valid = conv_read_0_cmd_valid;
  assign asMem_reads_0_sync_port_cmd_payload = conv_read_0_cmd_payload;
  assign conv_read_0_rsp = asMem_reads_0_sync_port_rsp;
  assign asMem_reads_1_sync_port_rsp = asMem_ram_spinal_port2;
  assign asMem_reads_1_sync_port_cmd_valid = conv_read_1_cmd_valid;
  assign asMem_reads_1_sync_port_cmd_payload = conv_read_1_cmd_payload;
  assign conv_read_1_rsp = asMem_reads_1_sync_port_rsp;

endmodule

module StreamArbiter_4 (
  input  wire          io_inputs_0_valid,
  output wire          io_inputs_0_ready,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [0:0]    io_chosenOH,
  input  wire          clk,
  input  wire          reset
);

  wire       [1:0]    _zz__zz_maskProposal_0_2;
  wire       [1:0]    _zz__zz_maskProposal_0_2_1;
  wire       [0:0]    _zz__zz_maskProposal_0_2_2;
  wire       [0:0]    _zz_maskProposal_0_3;
  reg                 locked;
  wire                maskProposal_0;
  reg                 maskLocked_0;
  wire                maskRouted_0;
  wire       [0:0]    _zz_maskProposal_0;
  wire       [1:0]    _zz_maskProposal_0_1;
  wire       [1:0]    _zz_maskProposal_0_2;
  wire                io_output_fire;

  assign _zz__zz_maskProposal_0_2 = (_zz_maskProposal_0_1 - _zz__zz_maskProposal_0_2_1);
  assign _zz__zz_maskProposal_0_2_2 = maskLocked_0;
  assign _zz__zz_maskProposal_0_2_1 = {1'd0, _zz__zz_maskProposal_0_2_2};
  assign _zz_maskProposal_0_3 = (_zz_maskProposal_0_2[1 : 1] | _zz_maskProposal_0_2[0 : 0]);
  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign _zz_maskProposal_0 = io_inputs_0_valid;
  assign _zz_maskProposal_0_1 = {_zz_maskProposal_0,_zz_maskProposal_0};
  assign _zz_maskProposal_0_2 = (_zz_maskProposal_0_1 & (~ _zz__zz_maskProposal_0_2));
  assign maskProposal_0 = _zz_maskProposal_0_3[0];
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign io_output_valid = (io_inputs_0_valid && maskRouted_0);
  assign io_inputs_0_ready = ((1'b0 || maskRouted_0) && io_output_ready);
  assign io_chosenOH = maskRouted_0;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      locked <= 1'b0;
      maskLocked_0 <= 1'b1;
    end else begin
      if(io_output_valid) begin
        maskLocked_0 <= maskRouted_0;
      end
      if(io_output_valid) begin
        locked <= 1'b1;
      end
      if(io_output_fire) begin
        locked <= 1'b0;
      end
    end
  end


endmodule

module StreamArbiter_3 (
  input  wire          io_inputs_0_valid,
  output wire          io_inputs_0_ready,
  input  wire [38:0]   io_inputs_0_payload_address,
  input  wire [0:0]    io_inputs_0_payload_storageId,
  input  wire          io_inputs_0_payload_storageEnable,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [38:0]   io_output_payload_address,
  output wire [0:0]    io_output_payload_storageId,
  output wire          io_output_payload_storageEnable,
  output wire [0:0]    io_chosenOH,
  input  wire          clk,
  input  wire          reset
);

  wire       [1:0]    _zz__zz_maskProposal_0_2;
  wire       [1:0]    _zz__zz_maskProposal_0_2_1;
  wire       [0:0]    _zz__zz_maskProposal_0_2_2;
  wire       [0:0]    _zz_maskProposal_0_3;
  reg                 locked;
  wire                maskProposal_0;
  reg                 maskLocked_0;
  wire                maskRouted_0;
  wire       [0:0]    _zz_maskProposal_0;
  wire       [1:0]    _zz_maskProposal_0_1;
  wire       [1:0]    _zz_maskProposal_0_2;
  wire                io_output_fire;

  assign _zz__zz_maskProposal_0_2 = (_zz_maskProposal_0_1 - _zz__zz_maskProposal_0_2_1);
  assign _zz__zz_maskProposal_0_2_2 = maskLocked_0;
  assign _zz__zz_maskProposal_0_2_1 = {1'd0, _zz__zz_maskProposal_0_2_2};
  assign _zz_maskProposal_0_3 = (_zz_maskProposal_0_2[1 : 1] | _zz_maskProposal_0_2[0 : 0]);
  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign _zz_maskProposal_0 = io_inputs_0_valid;
  assign _zz_maskProposal_0_1 = {_zz_maskProposal_0,_zz_maskProposal_0};
  assign _zz_maskProposal_0_2 = (_zz_maskProposal_0_1 & (~ _zz__zz_maskProposal_0_2));
  assign maskProposal_0 = _zz_maskProposal_0_3[0];
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign io_output_valid = (io_inputs_0_valid && maskRouted_0);
  assign io_output_payload_address = io_inputs_0_payload_address;
  assign io_output_payload_storageId = io_inputs_0_payload_storageId;
  assign io_output_payload_storageEnable = io_inputs_0_payload_storageEnable;
  assign io_inputs_0_ready = ((1'b0 || maskRouted_0) && io_output_ready);
  assign io_chosenOH = maskRouted_0;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      locked <= 1'b0;
      maskLocked_0 <= 1'b1;
    end else begin
      if(io_output_valid) begin
        maskLocked_0 <= maskRouted_0;
      end
      if(io_output_valid) begin
        locked <= 1'b1;
      end
      if(io_output_fire) begin
        locked <= 1'b0;
      end
    end
  end


endmodule

module StreamArbiter_2 (
  input  wire          io_inputs_0_valid,
  output wire          io_inputs_0_ready,
  input  wire [38:0]   io_inputs_0_payload_pcOnLastSlice,
  input  wire [38:0]   io_inputs_0_payload_pcTarget,
  input  wire          io_inputs_0_payload_taken,
  input  wire          io_inputs_0_payload_isBranch,
  input  wire          io_inputs_0_payload_isPush,
  input  wire          io_inputs_0_payload_isPop,
  input  wire          io_inputs_0_payload_wasWrong,
  input  wire          io_inputs_0_payload_badPredictedTarget,
  input  wire [11:0]   io_inputs_0_payload_history,
  input  wire [15:0]   io_inputs_0_payload_uopId,
  input  wire [1:0]    io_inputs_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_0,
  input  wire [1:0]    io_inputs_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_1,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [38:0]   io_output_payload_pcOnLastSlice,
  output wire [38:0]   io_output_payload_pcTarget,
  output wire          io_output_payload_taken,
  output wire          io_output_payload_isBranch,
  output wire          io_output_payload_isPush,
  output wire          io_output_payload_isPop,
  output wire          io_output_payload_wasWrong,
  output wire          io_output_payload_badPredictedTarget,
  output wire [11:0]   io_output_payload_history,
  output wire [15:0]   io_output_payload_uopId,
  output wire [1:0]    io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_0,
  output wire [1:0]    io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_1,
  output wire [0:0]    io_chosenOH,
  input  wire          clk,
  input  wire          reset
);

  wire       [1:0]    _zz__zz_maskProposal_0_2;
  wire       [1:0]    _zz__zz_maskProposal_0_2_1;
  wire       [0:0]    _zz__zz_maskProposal_0_2_2;
  wire       [0:0]    _zz_maskProposal_0_3;
  wire                locked;
  wire                maskProposal_0;
  reg                 maskLocked_0;
  wire                maskRouted_0;
  wire       [0:0]    _zz_maskProposal_0;
  wire       [1:0]    _zz_maskProposal_0_1;
  wire       [1:0]    _zz_maskProposal_0_2;

  assign _zz__zz_maskProposal_0_2 = (_zz_maskProposal_0_1 - _zz__zz_maskProposal_0_2_1);
  assign _zz__zz_maskProposal_0_2_2 = maskLocked_0;
  assign _zz__zz_maskProposal_0_2_1 = {1'd0, _zz__zz_maskProposal_0_2_2};
  assign _zz_maskProposal_0_3 = (_zz_maskProposal_0_2[1 : 1] | _zz_maskProposal_0_2[0 : 0]);
  assign locked = 1'b0;
  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign _zz_maskProposal_0 = io_inputs_0_valid;
  assign _zz_maskProposal_0_1 = {_zz_maskProposal_0,_zz_maskProposal_0};
  assign _zz_maskProposal_0_2 = (_zz_maskProposal_0_1 & (~ _zz__zz_maskProposal_0_2));
  assign maskProposal_0 = _zz_maskProposal_0_3[0];
  assign io_output_valid = (io_inputs_0_valid && maskRouted_0);
  assign io_output_payload_pcOnLastSlice = io_inputs_0_payload_pcOnLastSlice;
  assign io_output_payload_pcTarget = io_inputs_0_payload_pcTarget;
  assign io_output_payload_taken = io_inputs_0_payload_taken;
  assign io_output_payload_isBranch = io_inputs_0_payload_isBranch;
  assign io_output_payload_isPush = io_inputs_0_payload_isPush;
  assign io_output_payload_isPop = io_inputs_0_payload_isPop;
  assign io_output_payload_wasWrong = io_inputs_0_payload_wasWrong;
  assign io_output_payload_badPredictedTarget = io_inputs_0_payload_badPredictedTarget;
  assign io_output_payload_history = io_inputs_0_payload_history;
  assign io_output_payload_uopId = io_inputs_0_payload_uopId;
  assign io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 = io_inputs_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  assign io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_1 = io_inputs_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  assign io_inputs_0_ready = ((1'b0 || maskRouted_0) && io_output_ready);
  assign io_chosenOH = maskRouted_0;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      maskLocked_0 <= 1'b1;
    end else begin
      if(io_output_valid) begin
        maskLocked_0 <= maskRouted_0;
      end
    end
  end


endmodule

module StreamArbiter_1 (
  input  wire          io_inputs_0_valid,
  output wire          io_inputs_0_ready,
  input  wire [2:0]    io_inputs_0_payload_op,
  input  wire [38:0]   io_inputs_0_payload_address,
  input  wire [1:0]    io_inputs_0_payload_size,
  input  wire          io_inputs_0_payload_load,
  input  wire          io_inputs_0_payload_store,
  input  wire          io_inputs_0_payload_atomic,
  input  wire          io_inputs_0_payload_clean,
  input  wire          io_inputs_0_payload_invalidate,
  input  wire [11:0]   io_inputs_0_payload_storeId,
  input  wire          io_inputs_1_valid,
  output wire          io_inputs_1_ready,
  input  wire [2:0]    io_inputs_1_payload_op,
  input  wire [38:0]   io_inputs_1_payload_address,
  input  wire [1:0]    io_inputs_1_payload_size,
  input  wire          io_inputs_1_payload_load,
  input  wire          io_inputs_1_payload_store,
  input  wire          io_inputs_1_payload_atomic,
  input  wire          io_inputs_1_payload_clean,
  input  wire          io_inputs_1_payload_invalidate,
  input  wire [11:0]   io_inputs_1_payload_storeId,
  input  wire          io_inputs_2_valid,
  output wire          io_inputs_2_ready,
  input  wire [2:0]    io_inputs_2_payload_op,
  input  wire [38:0]   io_inputs_2_payload_address,
  input  wire [1:0]    io_inputs_2_payload_size,
  input  wire          io_inputs_2_payload_load,
  input  wire          io_inputs_2_payload_store,
  input  wire          io_inputs_2_payload_atomic,
  input  wire          io_inputs_2_payload_clean,
  input  wire          io_inputs_2_payload_invalidate,
  input  wire [11:0]   io_inputs_2_payload_storeId,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [2:0]    io_output_payload_op,
  output wire [38:0]   io_output_payload_address,
  output wire [1:0]    io_output_payload_size,
  output wire          io_output_payload_load,
  output wire          io_output_payload_store,
  output wire          io_output_payload_atomic,
  output wire          io_output_payload_clean,
  output wire          io_output_payload_invalidate,
  output wire [11:0]   io_output_payload_storeId,
  output wire [1:0]    io_chosen,
  output wire [2:0]    io_chosenOH,
  input  wire          clk,
  input  wire          reset
);
  localparam LsuL1CmdOpcode_LSU = 3'd0;
  localparam LsuL1CmdOpcode_ACCESS_1 = 3'd1;
  localparam LsuL1CmdOpcode_STORE_BUFFER = 3'd2;
  localparam LsuL1CmdOpcode_FLUSH = 3'd3;
  localparam LsuL1CmdOpcode_PREFETCH = 3'd4;

  wire       [2:0]    _zz__zz_maskProposal_1_1;
  reg        [2:0]    _zz__zz_io_output_payload_op;
  reg        [38:0]   _zz_io_output_payload_address_1;
  reg        [1:0]    _zz_io_output_payload_size;
  reg                 _zz_io_output_payload_load;
  reg                 _zz_io_output_payload_store;
  reg                 _zz_io_output_payload_atomic;
  reg                 _zz_io_output_payload_clean;
  reg                 _zz_io_output_payload_invalidate;
  reg        [11:0]   _zz_io_output_payload_storeId;
  wire                locked;
  wire                maskProposal_0;
  wire                maskProposal_1;
  wire                maskProposal_2;
  reg                 maskLocked_0;
  reg                 maskLocked_1;
  reg                 maskLocked_2;
  wire                maskRouted_0;
  wire                maskRouted_1;
  wire                maskRouted_2;
  wire       [2:0]    _zz_maskProposal_1;
  wire       [2:0]    _zz_maskProposal_1_1;
  wire       [1:0]    _zz_io_output_payload_address;
  wire       [2:0]    _zz_io_output_payload_op;
  wire                _zz_io_chosen;
  wire                _zz_io_chosen_1;
  `ifndef SYNTHESIS
  reg [95:0] io_inputs_0_payload_op_string;
  reg [95:0] io_inputs_1_payload_op_string;
  reg [95:0] io_inputs_2_payload_op_string;
  reg [95:0] io_output_payload_op_string;
  reg [95:0] _zz_io_output_payload_op_string;
  `endif


  assign _zz__zz_maskProposal_1_1 = (_zz_maskProposal_1 - 3'b001);
  always @(*) begin
    case(_zz_io_output_payload_address)
      2'b00 : begin
        _zz__zz_io_output_payload_op = io_inputs_0_payload_op;
        _zz_io_output_payload_address_1 = io_inputs_0_payload_address;
        _zz_io_output_payload_size = io_inputs_0_payload_size;
        _zz_io_output_payload_load = io_inputs_0_payload_load;
        _zz_io_output_payload_store = io_inputs_0_payload_store;
        _zz_io_output_payload_atomic = io_inputs_0_payload_atomic;
        _zz_io_output_payload_clean = io_inputs_0_payload_clean;
        _zz_io_output_payload_invalidate = io_inputs_0_payload_invalidate;
        _zz_io_output_payload_storeId = io_inputs_0_payload_storeId;
      end
      2'b01 : begin
        _zz__zz_io_output_payload_op = io_inputs_1_payload_op;
        _zz_io_output_payload_address_1 = io_inputs_1_payload_address;
        _zz_io_output_payload_size = io_inputs_1_payload_size;
        _zz_io_output_payload_load = io_inputs_1_payload_load;
        _zz_io_output_payload_store = io_inputs_1_payload_store;
        _zz_io_output_payload_atomic = io_inputs_1_payload_atomic;
        _zz_io_output_payload_clean = io_inputs_1_payload_clean;
        _zz_io_output_payload_invalidate = io_inputs_1_payload_invalidate;
        _zz_io_output_payload_storeId = io_inputs_1_payload_storeId;
      end
      default : begin
        _zz__zz_io_output_payload_op = io_inputs_2_payload_op;
        _zz_io_output_payload_address_1 = io_inputs_2_payload_address;
        _zz_io_output_payload_size = io_inputs_2_payload_size;
        _zz_io_output_payload_load = io_inputs_2_payload_load;
        _zz_io_output_payload_store = io_inputs_2_payload_store;
        _zz_io_output_payload_atomic = io_inputs_2_payload_atomic;
        _zz_io_output_payload_clean = io_inputs_2_payload_clean;
        _zz_io_output_payload_invalidate = io_inputs_2_payload_invalidate;
        _zz_io_output_payload_storeId = io_inputs_2_payload_storeId;
      end
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_inputs_0_payload_op)
      LsuL1CmdOpcode_LSU : io_inputs_0_payload_op_string = "LSU         ";
      LsuL1CmdOpcode_ACCESS_1 : io_inputs_0_payload_op_string = "ACCESS_1    ";
      LsuL1CmdOpcode_STORE_BUFFER : io_inputs_0_payload_op_string = "STORE_BUFFER";
      LsuL1CmdOpcode_FLUSH : io_inputs_0_payload_op_string = "FLUSH       ";
      LsuL1CmdOpcode_PREFETCH : io_inputs_0_payload_op_string = "PREFETCH    ";
      default : io_inputs_0_payload_op_string = "????????????";
    endcase
  end
  always @(*) begin
    case(io_inputs_1_payload_op)
      LsuL1CmdOpcode_LSU : io_inputs_1_payload_op_string = "LSU         ";
      LsuL1CmdOpcode_ACCESS_1 : io_inputs_1_payload_op_string = "ACCESS_1    ";
      LsuL1CmdOpcode_STORE_BUFFER : io_inputs_1_payload_op_string = "STORE_BUFFER";
      LsuL1CmdOpcode_FLUSH : io_inputs_1_payload_op_string = "FLUSH       ";
      LsuL1CmdOpcode_PREFETCH : io_inputs_1_payload_op_string = "PREFETCH    ";
      default : io_inputs_1_payload_op_string = "????????????";
    endcase
  end
  always @(*) begin
    case(io_inputs_2_payload_op)
      LsuL1CmdOpcode_LSU : io_inputs_2_payload_op_string = "LSU         ";
      LsuL1CmdOpcode_ACCESS_1 : io_inputs_2_payload_op_string = "ACCESS_1    ";
      LsuL1CmdOpcode_STORE_BUFFER : io_inputs_2_payload_op_string = "STORE_BUFFER";
      LsuL1CmdOpcode_FLUSH : io_inputs_2_payload_op_string = "FLUSH       ";
      LsuL1CmdOpcode_PREFETCH : io_inputs_2_payload_op_string = "PREFETCH    ";
      default : io_inputs_2_payload_op_string = "????????????";
    endcase
  end
  always @(*) begin
    case(io_output_payload_op)
      LsuL1CmdOpcode_LSU : io_output_payload_op_string = "LSU         ";
      LsuL1CmdOpcode_ACCESS_1 : io_output_payload_op_string = "ACCESS_1    ";
      LsuL1CmdOpcode_STORE_BUFFER : io_output_payload_op_string = "STORE_BUFFER";
      LsuL1CmdOpcode_FLUSH : io_output_payload_op_string = "FLUSH       ";
      LsuL1CmdOpcode_PREFETCH : io_output_payload_op_string = "PREFETCH    ";
      default : io_output_payload_op_string = "????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_output_payload_op)
      LsuL1CmdOpcode_LSU : _zz_io_output_payload_op_string = "LSU         ";
      LsuL1CmdOpcode_ACCESS_1 : _zz_io_output_payload_op_string = "ACCESS_1    ";
      LsuL1CmdOpcode_STORE_BUFFER : _zz_io_output_payload_op_string = "STORE_BUFFER";
      LsuL1CmdOpcode_FLUSH : _zz_io_output_payload_op_string = "FLUSH       ";
      LsuL1CmdOpcode_PREFETCH : _zz_io_output_payload_op_string = "PREFETCH    ";
      default : _zz_io_output_payload_op_string = "????????????";
    endcase
  end
  `endif

  assign locked = 1'b0;
  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskRouted_1 = (locked ? maskLocked_1 : maskProposal_1);
  assign maskRouted_2 = (locked ? maskLocked_2 : maskProposal_2);
  assign _zz_maskProposal_1 = {io_inputs_2_valid,{io_inputs_1_valid,io_inputs_0_valid}};
  assign _zz_maskProposal_1_1 = (_zz_maskProposal_1 & (~ _zz__zz_maskProposal_1_1));
  assign maskProposal_0 = io_inputs_0_valid;
  assign maskProposal_1 = _zz_maskProposal_1_1[1];
  assign maskProposal_2 = _zz_maskProposal_1_1[2];
  assign io_output_valid = (((io_inputs_0_valid && maskRouted_0) || (io_inputs_1_valid && maskRouted_1)) || (io_inputs_2_valid && maskRouted_2));
  assign _zz_io_output_payload_address = {maskRouted_2,maskRouted_1};
  assign _zz_io_output_payload_op = _zz__zz_io_output_payload_op;
  assign io_output_payload_op = _zz_io_output_payload_op;
  assign io_output_payload_address = _zz_io_output_payload_address_1;
  assign io_output_payload_size = _zz_io_output_payload_size;
  assign io_output_payload_load = _zz_io_output_payload_load;
  assign io_output_payload_store = _zz_io_output_payload_store;
  assign io_output_payload_atomic = _zz_io_output_payload_atomic;
  assign io_output_payload_clean = _zz_io_output_payload_clean;
  assign io_output_payload_invalidate = _zz_io_output_payload_invalidate;
  assign io_output_payload_storeId = _zz_io_output_payload_storeId;
  assign io_inputs_0_ready = ((1'b0 || maskRouted_0) && io_output_ready);
  assign io_inputs_1_ready = ((1'b0 || maskRouted_1) && io_output_ready);
  assign io_inputs_2_ready = ((1'b0 || maskRouted_2) && io_output_ready);
  assign io_chosenOH = {maskRouted_2,{maskRouted_1,maskRouted_0}};
  assign _zz_io_chosen = io_chosenOH[1];
  assign _zz_io_chosen_1 = io_chosenOH[2];
  assign io_chosen = {_zz_io_chosen_1,_zz_io_chosen};
  always @(posedge clk) begin
    if(io_output_valid) begin
      maskLocked_0 <= maskRouted_0;
      maskLocked_1 <= maskRouted_1;
      maskLocked_2 <= maskRouted_2;
    end
  end


endmodule

module StreamArbiter (
  input  wire          io_inputs_0_valid,
  output wire          io_inputs_0_ready,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [0:0]    io_chosenOH,
  input  wire          clk,
  input  wire          reset
);

  reg                 locked;
  wire                maskProposal_0;
  reg                 maskLocked_0;
  wire                maskRouted_0;
  wire                io_output_fire;

  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskProposal_0 = io_inputs_0_valid;
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign io_output_valid = (io_inputs_0_valid && maskRouted_0);
  assign io_inputs_0_ready = ((1'b0 || maskRouted_0) && io_output_ready);
  assign io_chosenOH = maskRouted_0;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      locked <= 1'b0;
    end else begin
      if(io_output_valid) begin
        locked <= 1'b1;
      end
      if(io_output_fire) begin
        locked <= 1'b0;
      end
    end
  end

  always @(posedge clk) begin
    if(io_output_valid) begin
      maskLocked_0 <= maskRouted_0;
    end
  end


endmodule

module DivRadix (
  input  wire          io_flush,
  input  wire          io_cmd_valid,
  output wire          io_cmd_ready,
  input  wire [63:0]   io_cmd_payload_a,
  input  wire [63:0]   io_cmd_payload_b,
  input  wire          io_cmd_payload_normalized,
  input  wire [5:0]    io_cmd_payload_iterations,
  output wire          io_rsp_valid,
  input  wire          io_rsp_ready,
  output wire [63:0]   io_rsp_payload_result,
  output wire [63:0]   io_rsp_payload_remain,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz_shifter_1;
  wire       [31:0]   _zz_shifter_2;
  wire       [47:0]   _zz_shifter_3;
  wire       [62:0]   _zz_shifter_4;
  reg        [5:0]    counter;
  reg                 busy;
  wire                io_rsp_fire;
  reg                 done;
  wire                when_DivRadix_l45;
  reg        [63:0]   shifter;
  reg        [63:0]   numerator;
  reg        [63:0]   result;
  reg        [64:0]   div1;
  reg        [64:0]   div3;
  wire       [64:0]   div2;
  wire       [64:0]   shifted;
  wire       [65:0]   sub1;
  wire                when_DivRadix_l64;
  reg        [64:0]   _zz_shifter;
  wire                when_DivRadix_l68;
  wire                slicesZero_0;
  wire                slicesZero_1;
  wire                slicesZero_2;
  wire       [2:0]    shiftSel;
  wire       [3:0]    _zz_sel;
  wire                _zz_sel_1;
  wire                _zz_sel_2;
  wire                _zz_sel_3;
  reg        [3:0]    _zz_sel_4;
  wire       [3:0]    _zz_sel_5;
  wire                _zz_sel_6;
  wire                _zz_sel_7;
  wire                _zz_sel_8;
  wire       [1:0]    sel;
  reg                 wasBusy;
  wire                when_DivRadix_l93;

  assign _zz_shifter_1 = io_cmd_payload_a[63 : 48];
  assign _zz_shifter_2 = io_cmd_payload_a[63 : 32];
  assign _zz_shifter_3 = io_cmd_payload_a[63 : 16];
  assign _zz_shifter_4 = io_cmd_payload_a[63 : 1];
  assign io_rsp_fire = (io_rsp_valid && io_rsp_ready);
  assign when_DivRadix_l45 = (busy && (counter == 6'h3f));
  assign div2 = (div1 <<< 1);
  assign shifted = {shifter,numerator[63 : 63]};
  assign sub1 = ({1'b0,shifted} - {1'b0,div1});
  assign io_rsp_valid = done;
  assign io_rsp_payload_result = result;
  assign io_rsp_payload_remain = shifter;
  assign io_cmd_ready = (! busy);
  assign when_DivRadix_l64 = (! done);
  always @(*) begin
    _zz_shifter = shifted;
    if(when_DivRadix_l68) begin
      _zz_shifter = sub1[64:0];
    end
  end

  assign when_DivRadix_l68 = (! sub1[65]);
  assign slicesZero_0 = (io_cmd_payload_a[31 : 16] == 16'h0);
  assign slicesZero_1 = (io_cmd_payload_a[47 : 32] == 16'h0);
  assign slicesZero_2 = (io_cmd_payload_a[63 : 48] == 16'h0);
  assign shiftSel = {(&slicesZero_2),{(&{slicesZero_2,slicesZero_1}),(&{slicesZero_2,{slicesZero_1,slicesZero_0}})}};
  assign _zz_sel = {1'b1,shiftSel};
  assign _zz_sel_1 = _zz_sel[0];
  assign _zz_sel_2 = _zz_sel[1];
  assign _zz_sel_3 = _zz_sel[2];
  always @(*) begin
    _zz_sel_4[0] = (_zz_sel_1 && (! 1'b0));
    _zz_sel_4[1] = (_zz_sel_2 && (! _zz_sel_1));
    _zz_sel_4[2] = (_zz_sel_3 && (! (|{_zz_sel_2,_zz_sel_1})));
    _zz_sel_4[3] = (_zz_sel[3] && (! (|{_zz_sel_3,{_zz_sel_2,_zz_sel_1}})));
  end

  assign _zz_sel_5 = _zz_sel_4;
  assign _zz_sel_6 = _zz_sel_5[3];
  assign _zz_sel_7 = (_zz_sel_5[1] || _zz_sel_6);
  assign _zz_sel_8 = (_zz_sel_5[2] || _zz_sel_6);
  assign sel = {_zz_sel_8,_zz_sel_7};
  assign when_DivRadix_l93 = (! busy);
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      busy <= 1'b0;
      done <= 1'b0;
      wasBusy <= 1'b0;
    end else begin
      if(io_rsp_fire) begin
        busy <= 1'b0;
      end
      if(when_DivRadix_l45) begin
        done <= 1'b1;
      end
      if(io_rsp_fire) begin
        done <= 1'b0;
      end
      wasBusy <= busy;
      if(when_DivRadix_l93) begin
        busy <= io_cmd_valid;
      end
      if(io_flush) begin
        done <= 1'b0;
        busy <= 1'b0;
      end
    end
  end

  always @(posedge clk) begin
    if(when_DivRadix_l64) begin
      counter <= (counter + 6'h01);
      result <= (result <<< 1);
      if(when_DivRadix_l68) begin
        result[0 : 0] <= 1'b1;
      end
      shifter <= _zz_shifter[63:0];
      numerator <= (numerator <<< 1);
    end
    if(when_DivRadix_l93) begin
      div1 <= {1'd0, io_cmd_payload_b};
      result <= ((io_cmd_payload_b == 64'h0) ? 64'hffffffffffffffff : 64'h0);
      case(sel)
        2'b11 : begin
          counter <= 6'h0;
          shifter <= 64'h0;
          numerator <= (io_cmd_payload_a <<< 0);
        end
        2'b10 : begin
          counter <= 6'h10;
          shifter <= {48'd0, _zz_shifter_1};
          numerator <= (io_cmd_payload_a <<< 16);
        end
        2'b01 : begin
          counter <= 6'h20;
          shifter <= {32'd0, _zz_shifter_2};
          numerator <= (io_cmd_payload_a <<< 32);
        end
        default : begin
          counter <= 6'h30;
          shifter <= {16'd0, _zz_shifter_3};
          numerator <= (io_cmd_payload_a <<< 48);
        end
      endcase
      if(io_cmd_payload_normalized) begin
        counter <= (6'h3f - io_cmd_payload_iterations);
        shifter <= {1'd0, _zz_shifter_4};
        numerator <= (io_cmd_payload_a <<< 63);
      end
    end
  end


endmodule
